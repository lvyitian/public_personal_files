module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_23), .en(wire_61), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_65), .in(arch_input_value), .out(wire_55));
  TC_Program8_4 # (.UUID(64'd4489305393227859486 ^ UUID), .DEFAULT_FILE_NAME("Program8_4_3E4D37784397861E.w8.bin"), .ARG_SIG("Program8_4_3E4D37784397861E=%s")) Program8_4_2 (.clk(clk), .rst(rst), .address(wire_2), .out0(wire_3), .out1(wire_1), .out2(wire_5), .out3(wire_48));
  TC_Counter # (.UUID(64'd1175999672554394000 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_3 (.clk(clk), .rst(rst), .save(wire_57), .in(wire_23), .out(wire_2));
  TC_Splitter8 # (.UUID(64'd3496280010280654809 ^ UUID)) Splitter8_4 (.in(wire_34), .out0(wire_64), .out1(wire_54), .out2(wire_58), .out3(wire_59), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1350359362790102949 ^ UUID)) Splitter8_5 (.in(wire_41), .out0(wire_11), .out1(wire_18), .out2(wire_60), .out3(wire_78), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3688384451292696869 ^ UUID)) Splitter8_6 (.in(wire_62), .out0(wire_66), .out1(wire_24), .out2(wire_26), .out3(wire_8), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3357720912797461292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_0), .in(wire_2), .out());
  TC_Maker8 # (.UUID(64'd2922775923237819214 ^ UUID)) Maker8_8 (.in0(wire_74), .in1(wire_79), .in2(wire_83), .in3(wire_40), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_36));
  TC_Splitter8 # (.UUID(64'd4136660363423911410 ^ UUID)) Splitter8_9 (.in(wire_3), .out0(wire_74), .out1(wire_79), .out2(wire_83), .out3(wire_40), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd4550958897663313502 ^ UUID)) Splitter8_10 (.in(wire_3), .out0(wire_77), .out1(wire_51), .out2(wire_30), .out3(wire_33), .out4(wire_56), .out5(wire_28), .out6(wire_69), .out7(wire_17));
  TC_Maker8 # (.UUID(64'd3153840370766490713 ^ UUID)) Maker8_11 (.in0(wire_77), .in1(wire_51), .in2(wire_30), .in3(wire_33), .in4(wire_56), .in5(wire_28), .in6(wire_69), .in7(wire_17), .out(wire_70));
  TC_Constant # (.UUID(64'd4029987529778329422 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out(wire_22));
  TC_Constant # (.UUID(64'd47372170638122597 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_81));
  TC_Constant # (.UUID(64'd3010400910295959985 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_7));
  TC_Constant # (.UUID(64'd1353887318054096472 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out(wire_71));
  TC_Constant # (.UUID(64'd4461919415197064488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_4));
  TC_Constant # (.UUID(64'd2551986311311524963 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out(wire_14));
  TC_Switch # (.UUID(64'd201407107924193690 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_45), .in(wire_21), .out(wire_27_0));
  TC_Switch # (.UUID(64'd3784926049681585699 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_47), .in(wire_21), .out(wire_9_1));
  TC_Switch # (.UUID(64'd3418942253385023549 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_15), .in(wire_38), .out(wire_27_2));
  TC_Switch # (.UUID(64'd3104771108315787100 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_32), .in(wire_38), .out(wire_9_0));
  TC_Switch # (.UUID(64'd494263610589549334 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_46), .in(wire_50), .out(wire_27_6));
  TC_Switch # (.UUID(64'd4455028313033582898 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_35), .in(wire_50), .out(wire_9_2));
  TC_Switch # (.UUID(64'd977062972681925203 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_68), .in(wire_37), .out(wire_27_3));
  TC_Switch # (.UUID(64'd2935373336597064260 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_25), .in(wire_37), .out(wire_9_4));
  TC_Switch # (.UUID(64'd2595310988575568445 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_19), .in(wire_43), .out(wire_27_5));
  TC_Switch # (.UUID(64'd3649926646471230167 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_63), .in(wire_43), .out(wire_9_3));
  TC_Switch # (.UUID(64'd115863760055946247 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_31), .in(wire_52), .out(wire_27_7));
  TC_Switch # (.UUID(64'd459043271910661458 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_73), .in(wire_52), .out(wire_9_5));
  TC_Switch # (.UUID(64'd4275937720180353902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_80), .in(wire_2), .out());
  TC_Switch # (.UUID(64'd2718446434835356700 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_13), .in(wire_55), .out(wire_27_4));
  TC_Switch # (.UUID(64'd1811299859375739998 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_42), .in(wire_55), .out(wire_9_6));
  TC_Or # (.UUID(64'd117421755651659184 ^ UUID), .BIT_WIDTH(64'd1)) Or_33 (.in0(wire_13), .in1(wire_42), .out(wire_65));
  TC_Switch # (.UUID(64'd262409980643160938 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_12), .in(wire_5), .out(wire_9_7));
  TC_Switch # (.UUID(64'd2764614579549035605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_53), .in(wire_1), .out(wire_27_1));
  TC_Switch # (.UUID(64'd2974460371787013801 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_29), .in(wire_44), .out(wire_23_1));
  TC_Mux # (.UUID(64'd1769789085559769130 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_37 (.sel(wire_12), .in0(wire_5), .in1(wire_82), .out(wire_41));
  TC_Mux # (.UUID(64'd1404337327044278632 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_53), .in0(wire_1), .in1(wire_75), .out(wire_34));
  TC_Constant # (.UUID(64'd4387708643330744374 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_39 (.out(wire_75));
  TC_Constant # (.UUID(64'd2430039925245603401 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_40 (.out(wire_82));
  TC_Switch # (.UUID(64'd3877536405880520929 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_67), .in(wire_6), .out(wire_16));
  TC_Constant # (.UUID(64'd2430392602802046886 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_42 (.out(wire_72));
  TC_Mux # (.UUID(64'd1559488034901936773 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_43 (.sel(wire_16), .in0(wire_48), .in1(wire_72), .out(wire_62));
  TC_Switch # (.UUID(64'd3981948550050450551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_16), .in(wire_48), .out(wire_23_0));
  _4bit_Decoder # (.UUID(64'd188593635878702660 ^ UUID)) _4bit_Decoder_45 (.clk(clk), .rst(rst), .\1_1 (wire_64), .\2_1 (wire_54), .\4_1 (wire_58), .\8_1 (wire_59), .\7 (wire_13), .\11 (), .\3 (wire_68), .\15 (), .\6 (wire_0), .\8_2 (), .\5 (wire_31), .\9 (), .\10 (), .\4_2 (wire_19), .\12 (), .\13 (), .\14 (), .\2_2 (wire_46), .\1_2 (wire_15), .\0 (wire_45));
  _4bit_Decoder # (.UUID(64'd3657203059375966986 ^ UUID)) _4bit_Decoder_46 (.clk(clk), .rst(rst), .\1_1 (wire_11), .\2_1 (wire_18), .\4_1 (wire_60), .\8_1 (wire_78), .\7 (wire_42), .\11 (), .\3 (wire_25), .\15 (), .\6 (wire_80), .\8_2 (), .\5 (wire_73), .\9 (), .\10 (), .\4_2 (wire_63), .\12 (), .\13 (), .\14 (), .\2_2 (wire_35), .\1_2 (wire_32), .\0 (wire_47));
  _4bit_Decoder # (.UUID(64'd4526675728054865805 ^ UUID)) _4bit_Decoder_47 (.clk(clk), .rst(rst), .\1_1 (wire_66), .\2_1 (wire_24), .\4_1 (wire_26), .\8_1 (wire_8), .\7 (wire_61), .\11 (), .\3 (wire_49), .\15 (), .\6 (wire_57), .\8_2 (), .\5 (wire_39), .\9 (), .\10 (), .\4_2 (wire_76), .\12 (), .\13 (), .\14 (), .\2_2 (wire_84), .\1_2 (wire_20), .\0 (wire_10));
  RegisterPlus # (.UUID(64'd1898575026262245003 ^ UUID)) RegisterPlus_48 (.clk(clk), .rst(rst), .\�_____ (wire_22), .\�___________ (wire_23), .\�_____ (wire_10), .\�___________ (), .Output(wire_21));
  RegisterPlus # (.UUID(64'd201486149512558618 ^ UUID)) RegisterPlus_49 (.clk(clk), .rst(rst), .\�_____ (wire_81), .\�___________ (wire_23), .\�_____ (wire_20), .\�___________ (), .Output(wire_38));
  RegisterPlus # (.UUID(64'd4130910523704063521 ^ UUID)) RegisterPlus_50 (.clk(clk), .rst(rst), .\�_____ (wire_7), .\�___________ (wire_23), .\�_____ (wire_84), .\�___________ (), .Output(wire_50));
  RegisterPlus # (.UUID(64'd579904311903668382 ^ UUID)) RegisterPlus_51 (.clk(clk), .rst(rst), .\�_____ (wire_71), .\�___________ (wire_23), .\�_____ (wire_49), .\�___________ (), .Output(wire_37));
  RegisterPlus # (.UUID(64'd2026589517635316452 ^ UUID)) RegisterPlus_52 (.clk(clk), .rst(rst), .\�_____ (wire_4), .\�___________ (wire_23), .\�_____ (wire_76), .\�___________ (), .Output(wire_43));
  RegisterPlus # (.UUID(64'd1622410096212380183 ^ UUID)) RegisterPlus_53 (.clk(clk), .rst(rst), .\�_____ (wire_14), .\�___________ (wire_23), .\�_____ (wire_39), .\�___________ (), .Output(wire_52));
  LEG_ALU # (.UUID(64'd740631443788402157 ^ UUID)) LEG_ALU_54 (.clk(clk), .rst(rst), .\�_____ (wire_36), .\�______1 (wire_27), .\�______2 (wire_9), .Output(wire_44));
  LEG_DEC # (.UUID(64'd1666076388199409894 ^ UUID)) LEG_DEC_55 (.clk(clk), .rst(rst), .OPCODE(wire_70), .IMMEDIATE1(wire_53), .IMMEDIATE2(wire_12), .CALCULATION(wire_29), .JUMP(wire_67));
  LEG_COND # (.UUID(64'd999600516743479399 ^ UUID)) LEG_COND_56 (.clk(clk), .rst(rst), .ARG1(wire_27), .ARG2(wire_9), .\�_____ (wire_3), .Output(wire_6));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_9_0;
  wire [7:0] wire_9_1;
  wire [7:0] wire_9_2;
  wire [7:0] wire_9_3;
  wire [7:0] wire_9_4;
  wire [7:0] wire_9_5;
  wire [7:0] wire_9_6;
  wire [7:0] wire_9_7;
  assign wire_9 = wire_9_0|wire_9_1|wire_9_2|wire_9_3|wire_9_4|wire_9_5|wire_9_6|wire_9_7;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_23_0;
  wire [7:0] wire_23_1;
  assign wire_23 = wire_23_0|wire_23_1;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_27_0;
  wire [7:0] wire_27_1;
  wire [7:0] wire_27_2;
  wire [7:0] wire_27_3;
  wire [7:0] wire_27_4;
  wire [7:0] wire_27_5;
  wire [7:0] wire_27_6;
  wire [7:0] wire_27_7;
  assign wire_27 = wire_27_0|wire_27_1|wire_27_2|wire_27_3|wire_27_4|wire_27_5|wire_27_6|wire_27_7;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  assign arch_output_enable = wire_61;
  wire [7:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  assign arch_input_enable = wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [7:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [7:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;

endmodule
