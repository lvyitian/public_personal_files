module LEG_COND (clk, rst, ARG1, ARG2, \�_____ , Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] ARG1;
  input  wire [7:0] ARG2;
  input  wire [7:0] \�_____ ;
  output  wire [0:0] Output;

  TC_Equal # (.UUID(64'd469022450449281397 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_0 (.in0(wire_4), .in1(wire_32), .out(wire_27));
  TC_Constant # (.UUID(64'd2051448023974927123 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h20)) Constant8_1 (.out(wire_32));
  TC_Equal # (.UUID(64'd302087503831493541 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_2 (.in0(wire_4), .in1(wire_30), .out(wire_18));
  TC_Constant # (.UUID(64'd4542222613295176889 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h21)) Constant8_3 (.out(wire_30));
  TC_Equal # (.UUID(64'd3977699302148921626 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_4 (.in0(wire_4), .in1(wire_24), .out(wire_21));
  TC_Constant # (.UUID(64'd2314937324333883295 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h22)) Constant8_5 (.out(wire_24));
  TC_Equal # (.UUID(64'd2598179579939704549 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_6 (.in0(wire_4), .in1(wire_14), .out(wire_38));
  TC_Constant # (.UUID(64'd2619140119885518802 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h23)) Constant8_7 (.out(wire_14));
  TC_Equal # (.UUID(64'd1016355148453492596 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_8 (.in0(wire_4), .in1(wire_22), .out(wire_29));
  TC_Constant # (.UUID(64'd1550705849817143486 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h24)) Constant8_9 (.out(wire_22));
  TC_Equal # (.UUID(64'd1602625343120996724 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_10 (.in0(wire_4), .in1(wire_13), .out(wire_15));
  TC_Constant # (.UUID(64'd2222307270319111175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h25)) Constant8_11 (.out(wire_13));
  TC_Not # (.UUID(64'd2244182005895984404 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_11), .out(wire_8));
  TC_Equal # (.UUID(64'd168532653866922664 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_13 (.in0(wire_9), .in1(wire_7), .out(wire_11));
  TC_Switch # (.UUID(64'd859839441511864255 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_27), .in(wire_11), .out(wire_2_5));
  TC_Switch # (.UUID(64'd3687602544865986092 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_15 (.en(wire_18), .in(wire_8), .out(wire_2_8));
  TC_LessU # (.UUID(64'd2837489368470343284 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_16 (.in0(wire_9), .in1(wire_7), .out(wire_3));
  TC_Switch # (.UUID(64'd114564404545293814 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_21), .in(wire_3), .out(wire_2_7));
  TC_Switch # (.UUID(64'd3233876504730006742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_38), .in(wire_40), .out(wire_2_4));
  TC_Or # (.UUID(64'd1752390656836275508 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_3), .in1(wire_11), .out(wire_40));
  TC_Switch # (.UUID(64'd1313143816079393951 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_20 (.en(wire_15), .in(wire_0), .out(wire_2_9));
  TC_Not # (.UUID(64'd1225463839904331438 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_3), .out(wire_0));
  TC_Switch # (.UUID(64'd3591175240098488323 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_29), .in(wire_34), .out(wire_2_6));
  TC_And # (.UUID(64'd2923998825401666618 ^ UUID), .BIT_WIDTH(64'd1)) And_23 (.in0(wire_8), .in1(wire_0), .out(wire_34));
  TC_Maker8 # (.UUID(64'd4350048876850400171 ^ UUID)) Maker8_24 (.in0(wire_19), .in1(wire_16), .in2(wire_35), .in3(wire_36), .in4(wire_5), .in5(wire_31), .in6(1'd0), .in7(1'd0), .out(wire_4));
  TC_Splitter8 # (.UUID(64'd3964202440971776894 ^ UUID)) Splitter8_25 (.in(wire_33), .out0(wire_19), .out1(wire_16), .out2(wire_35), .out3(wire_36), .out4(wire_5), .out5(wire_31), .out6(), .out7());
  TC_Equal # (.UUID(64'd1260754848101083012 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_26 (.in0(wire_4), .in1(wire_10), .out(wire_17));
  TC_Constant # (.UUID(64'd980951910217902543 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h26)) Constant8_27 (.out(wire_10));
  TC_Constant # (.UUID(64'd2997422239060942000 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h27)) Constant8_28 (.out(wire_1));
  TC_Equal # (.UUID(64'd899453443110480878 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_29 (.in0(wire_4), .in1(wire_1), .out(wire_25));
  TC_Constant # (.UUID(64'd2927950784883307602 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h28)) Constant8_30 (.out(wire_23));
  TC_Equal # (.UUID(64'd241406386753268791 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_31 (.in0(wire_4), .in1(wire_23), .out(wire_39));
  TC_Constant # (.UUID(64'd4145911819613088554 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h29)) Constant8_32 (.out(wire_26));
  TC_Equal # (.UUID(64'd2085230340721355945 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_33 (.in0(wire_4), .in1(wire_26), .out(wire_28));
  TC_Switch # (.UUID(64'd3789360908499522547 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_17), .in(wire_6), .out(wire_2_3));
  TC_Switch # (.UUID(64'd257917569845715035 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_35 (.en(wire_25), .in(wire_20), .out(wire_2_2));
  TC_Switch # (.UUID(64'd2095736601766047070 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_39), .in(wire_37), .out(wire_2_0));
  TC_Switch # (.UUID(64'd3716747265466847797 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_37 (.en(wire_28), .in(wire_12), .out(wire_2_1));
  TC_LessI # (.UUID(64'd1385355206190587062 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_38 (.in0(wire_9), .in1(wire_7), .out(wire_6));
  TC_Or # (.UUID(64'd3012749455494048092 ^ UUID), .BIT_WIDTH(64'd1)) Or_39 (.in0(wire_6), .in1(wire_11), .out(wire_20));
  TC_Not # (.UUID(64'd2249480345734393481 ^ UUID), .BIT_WIDTH(64'd1)) Not_40 (.in(wire_6), .out(wire_12));
  TC_And # (.UUID(64'd2947011798661445761 ^ UUID), .BIT_WIDTH(64'd1)) And_41 (.in0(wire_8), .in1(wire_12), .out(wire_37));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_2_0;
  wire [0:0] wire_2_1;
  wire [0:0] wire_2_2;
  wire [0:0] wire_2_3;
  wire [0:0] wire_2_4;
  wire [0:0] wire_2_5;
  wire [0:0] wire_2_6;
  wire [0:0] wire_2_7;
  wire [0:0] wire_2_8;
  wire [0:0] wire_2_9;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8|wire_2_9;
  assign Output = wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = ARG2;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  assign wire_9 = ARG1;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_33;
  assign wire_33 = \�_____ ;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;

endmodule
