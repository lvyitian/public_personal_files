module COND (clk, rst, \�_____ , \�______1 , \�______2 );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] \�_____ ;
  input  wire [7:0] \�______1 ;
  output  wire [0:0] \�______2 ;

  TC_Decoder3 # (.UUID(64'd2925115600376390304 ^ UUID)) Decoder3_0 (.dis(1'd0), .sel0(wire_43), .sel1(wire_22), .sel2(wire_0), .out0(), .out1(wire_20), .out2(wire_13), .out3(wire_4), .out4(wire_39), .out5(wire_29), .out6(wire_34), .out7(wire_27));
  TC_Splitter8 # (.UUID(64'd3470519188273703912 ^ UUID)) Splitter8_1 (.in(wire_25), .out0(wire_43), .out1(wire_22), .out2(wire_0), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd4334758234279334509 ^ UUID)) Splitter8_2 (.in(wire_23), .out0(wire_14), .out1(wire_31), .out2(wire_44), .out3(wire_7), .out4(wire_18), .out5(wire_6), .out6(wire_9), .out7(wire_21));
  TC_Not # (.UUID(64'd3356655775406523277 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_14), .out(wire_17));
  TC_Not # (.UUID(64'd3372003852346323509 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_31), .out(wire_37));
  TC_Not # (.UUID(64'd4300359231852631695 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_44), .out(wire_24));
  TC_Not # (.UUID(64'd4274228112083492922 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_7), .out(wire_40));
  TC_Not # (.UUID(64'd2902193455854584740 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_18), .out(wire_3));
  TC_Not # (.UUID(64'd228192272609183863 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_6), .out(wire_15));
  TC_Not # (.UUID(64'd798670888936031036 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_9), .out(wire_16));
  TC_Not # (.UUID(64'd1999972821766259893 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_21), .out(wire_28));
  TC_And3 # (.UUID(64'd2059677990304844505 ^ UUID), .BIT_WIDTH(64'd1)) And3_11 (.in0(wire_17), .in1(wire_37), .in2(wire_24), .out(wire_38));
  TC_And3 # (.UUID(64'd948522879768405750 ^ UUID), .BIT_WIDTH(64'd1)) And3_12 (.in0(wire_38), .in1(wire_40), .in2(wire_3), .out(wire_35));
  TC_And3 # (.UUID(64'd4372362206184088052 ^ UUID), .BIT_WIDTH(64'd1)) And3_13 (.in0(wire_35), .in1(wire_15), .in2(wire_16), .out(wire_5));
  TC_And # (.UUID(64'd3123548669855028618 ^ UUID), .BIT_WIDTH(64'd1)) And_14 (.in0(wire_5), .in1(wire_28), .out(wire_10));
  TC_Switch # (.UUID(64'd634679830248559241 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_15 (.en(wire_11), .in(wire_21), .out(wire_36));
  TC_Switch # (.UUID(64'd2795670288739424508 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_16 (.en(wire_19), .in(wire_10), .out(wire_8));
  TC_Or3 # (.UUID(64'd2306917535285242489 ^ UUID), .BIT_WIDTH(64'd1)) Or3_17 (.in0(wire_20), .in1(wire_4), .in2(wire_34), .out(wire_19));
  TC_Or # (.UUID(64'd3746409483646556895 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_13), .in1(wire_4), .out(wire_11));
  TC_Or3 # (.UUID(64'd3648234591776454774 ^ UUID), .BIT_WIDTH(64'd1)) Or3_19 (.in0(wire_8), .in1(wire_36), .in2(wire_39), .out(wire_42));
  TC_Switch # (.UUID(64'd4059939730348919149 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_20 (.en(wire_29), .in(wire_1), .out(wire_2));
  TC_Or3 # (.UUID(64'd1654113391022042074 ^ UUID), .BIT_WIDTH(64'd1)) Or3_21 (.in0(wire_42), .in1(wire_2), .in2(wire_26), .out(wire_32));
  TC_Not # (.UUID(64'd144925859667489712 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_10), .out(wire_1));
  TC_Switch # (.UUID(64'd2403630434640686559 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_23 (.en(wire_33), .in(wire_12), .out(wire_26));
  TC_Or # (.UUID(64'd4070071511209401408 ^ UUID), .BIT_WIDTH(64'd1)) Or_24 (.in0(wire_34), .in1(wire_27), .out(wire_33));
  TC_Not # (.UUID(64'd4321257432484836311 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_21), .out(wire_30));
  TC_And # (.UUID(64'd1755950260431621294 ^ UUID), .BIT_WIDTH(64'd1)) And_26 (.in0(wire_30), .in1(wire_41), .out(wire_12));
  TC_Not # (.UUID(64'd946478276252201397 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_10), .out(wire_41));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  assign wire_23 = \�______1 ;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  assign wire_25 = \�_____ ;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  assign \�______2  = wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;

endmodule
