module Instructionz_Decoder (clk, rst, Input, Enabled, ALU, Control, Memory_Read, Fence, System, Error);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Input;
  input  wire [0:0] Enabled;
  output  wire [0:0] ALU;
  output  wire [0:0] Control;
  output  wire [0:0] Memory_Read;
  output  wire [0:0] Fence;
  output  wire [0:0] System;
  output  wire [0:0] Error;

  TC_Splitter32 # (.UUID(64'd3947739734663349922 ^ UUID)) Splitter32_0 (.in(wire_44), .out0(wire_7), .out1(), .out2(), .out3());
  TC_Splitter8 # (.UUID(64'd3117991262660878578 ^ UUID)) Splitter8_1 (.in(wire_7), .out0(wire_14), .out1(wire_16), .out2(wire_10), .out3(wire_1), .out4(wire_11), .out5(wire_22), .out6(wire_4), .out7());
  TC_And3 # (.UUID(64'd980466729639594772 ^ UUID), .BIT_WIDTH(64'd1)) And3_2 (.in0(wire_13), .in1(wire_22), .in2(wire_4), .out(wire_9));
  TC_Not # (.UUID(64'd2340154427682436773 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_11), .out(wire_13));
  TC_Nand # (.UUID(64'd1801162032929421007 ^ UUID), .BIT_WIDTH(64'd1)) Nand_4 (.in0(wire_14), .in1(wire_16), .out(wire_33));
  TC_Not # (.UUID(64'd2210352776962588522 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_4), .out(wire_25));
  TC_Not # (.UUID(64'd4310025696028194660 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_1), .out(wire_17));
  TC_And # (.UUID(64'd149724151827786004 ^ UUID), .BIT_WIDTH(64'd1)) And_7 (.in0(wire_19), .in1(wire_34), .out(wire_8));
  TC_And # (.UUID(64'd190446292339745544 ^ UUID), .BIT_WIDTH(64'd1)) And_8 (.in0(wire_15), .in1(wire_43), .out(wire_19));
  TC_Not # (.UUID(64'd3498325639852527168 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_4), .out(wire_35));
  TC_Not # (.UUID(64'd1455884858090119196 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_11), .out(wire_23));
  TC_Not # (.UUID(64'd2087933824073351986 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_1), .out(wire_43));
  TC_Not # (.UUID(64'd3661043119746078253 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_10), .out(wire_15));
  TC_And3 # (.UUID(64'd3692189082489085542 ^ UUID), .BIT_WIDTH(64'd1)) And3_13 (.in0(wire_26), .in1(wire_32), .in2(wire_41), .out(wire_37));
  TC_And # (.UUID(64'd3259121963457519506 ^ UUID), .BIT_WIDTH(64'd1)) And_14 (.in0(wire_10), .in1(wire_1), .out(wire_27));
  TC_And # (.UUID(64'd4071735716691435052 ^ UUID), .BIT_WIDTH(64'd1)) And_15 (.in0(wire_27), .in1(wire_37), .out(wire_6));
  TC_Not # (.UUID(64'd4420977415501974783 ^ UUID), .BIT_WIDTH(64'd1)) Not_16 (.in(wire_4), .out(wire_41));
  TC_Not # (.UUID(64'd3617292458837153491 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_22), .out(wire_32));
  TC_Not # (.UUID(64'd129744789343158879 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_11), .out(wire_26));
  TC_And3 # (.UUID(64'd4085345558270935283 ^ UUID), .BIT_WIDTH(64'd1)) And3_19 (.in0(wire_11), .in1(wire_22), .in2(wire_4), .out(wire_21));
  TC_And # (.UUID(64'd4072668974764630127 ^ UUID), .BIT_WIDTH(64'd1)) And_20 (.in0(wire_31), .in1(wire_20), .out(wire_28));
  TC_And # (.UUID(64'd2066749772917604869 ^ UUID), .BIT_WIDTH(64'd1)) And_21 (.in0(wire_28), .in1(wire_21), .out(wire_0));
  TC_Not # (.UUID(64'd4546996868130193819 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_1), .out(wire_20));
  TC_Not # (.UUID(64'd810264584082682700 ^ UUID), .BIT_WIDTH(64'd1)) Not_23 (.in(wire_10), .out(wire_31));
  TC_And3 # (.UUID(64'd2073327864954767054 ^ UUID), .BIT_WIDTH(64'd1)) And3_24 (.in0(wire_17), .in1(wire_11), .in2(wire_25), .out(wire_3));
  TC_Or3 # (.UUID(64'd3971525562417407934 ^ UUID), .BIT_WIDTH(64'd1)) Or3_25 (.in0(wire_9), .in1(wire_3), .in2(wire_8), .out(wire_24));
  TC_Or3 # (.UUID(64'd1416107883033528113 ^ UUID), .BIT_WIDTH(64'd1)) Or3_26 (.in0(wire_6), .in1(wire_0), .in2(1'd0), .out(wire_30));
  TC_Or # (.UUID(64'd4152805452209084740 ^ UUID), .BIT_WIDTH(64'd1)) Or_27 (.in0(wire_24), .in1(wire_30), .out(wire_42));
  TC_Not # (.UUID(64'd1184562550084866268 ^ UUID), .BIT_WIDTH(64'd1)) Not_28 (.in(wire_42), .out(wire_18));
  TC_Or # (.UUID(64'd4565495870725328242 ^ UUID), .BIT_WIDTH(64'd1)) Or_29 (.in0(wire_33), .in1(wire_18), .out(wire_39));
  TC_And # (.UUID(64'd4121673666677999850 ^ UUID), .BIT_WIDTH(64'd1)) And_30 (.in0(wire_23), .in1(wire_35), .out(wire_34));
  TC_And # (.UUID(64'd2960061295601050077 ^ UUID), .BIT_WIDTH(64'd1)) And_31 (.in0(wire_5), .in1(wire_39), .out(wire_36));
  TC_Switch # (.UUID(64'd753838681169017655 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_32 (.en(wire_5), .in(wire_9), .out(wire_38));
  TC_Switch # (.UUID(64'd3995209055622036913 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_33 (.en(wire_5), .in(wire_3), .out(wire_2));
  TC_Switch # (.UUID(64'd2653717390643449863 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_5), .in(wire_8), .out(wire_29));
  TC_Switch # (.UUID(64'd228730318812683385 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_35 (.en(wire_5), .in(wire_6), .out(wire_12));
  TC_Switch # (.UUID(64'd3891761927353018975 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_5), .in(wire_0), .out(wire_40));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign ALU = wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  assign wire_5 = Enabled;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  assign Fence = wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  assign Memory_Read = wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  assign Error = wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  assign Control = wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  assign System = wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [31:0] wire_44;
  assign wire_44 = Input;

endmodule
