// Dummy implementation, does nothing
module TC_Console (clk, rst, offset);
    parameter UUID = 0;
    parameter NAME = "";
    input clk;
    input rst;
    input [31:0] offset;
endmodule
