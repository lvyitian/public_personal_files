module Displayz_Controller (clk, rst, Value, Enable, Address, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8, Output_9, Output_10, Output_11, Output_12, Output_13, Output_14, Output_15, Output_16, Output_17, Output_18, Output_19, Output_20, Output_21, Output_22, Output_23, Output_24);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Value;
  input  wire [0:0] Enable;
  input  wire [31:0] Address;
  output  wire [31:0] Output_1;
  output  wire [31:0] Output_2;
  output  wire [31:0] Output_3;
  output  wire [31:0] Output_4;
  output  wire [31:0] Output_5;
  output  wire [31:0] Output_6;
  output  wire [31:0] Output_7;
  output  wire [31:0] Output_8;
  output  wire [31:0] Output_9;
  output  wire [31:0] Output_10;
  output  wire [31:0] Output_11;
  output  wire [31:0] Output_12;
  output  wire [31:0] Output_13;
  output  wire [31:0] Output_14;
  output  wire [31:0] Output_15;
  output  wire [31:0] Output_16;
  output  wire [63:0] Output_17;
  output  wire [63:0] Output_18;
  output  wire [63:0] Output_19;
  output  wire [63:0] Output_20;
  output  wire [63:0] Output_21;
  output  wire [63:0] Output_22;
  output  wire [63:0] Output_23;
  output  wire [63:0] Output_24;

  TC_Mul # (.UUID(64'd998942097976894219 ^ UUID), .BIT_WIDTH(64'd32)) DivMod32_0 (.in0(wire_9), .in1(wire_77), .out0(wire_60), .out1(wire_43));
  TC_Constant # (.UUID(64'd1706953689208840521 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h60)) Constant32_1 (.out(wire_77));
  TC_Decoder3 # (.UUID(64'd3124819825474212326 ^ UUID)) Decoder3_2 (.dis(wire_22), .sel0(wire_42), .sel1(wire_23), .sel2(wire_12), .out0(wire_17), .out1(wire_98), .out2(wire_91), .out3(wire_86), .out4(wire_53), .out5(wire_7), .out6(wire_39), .out7(wire_56));
  TC_Splitter8 # (.UUID(64'd2689414568765749380 ^ UUID)) Splitter8_3 (.in(wire_31), .out0(wire_42), .out1(wire_23), .out2(wire_12), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2577865555952160451 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_75), .out(wire_22));
  TC_Constant # (.UUID(64'd2987616758561940336 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_5 (.out(wire_10));
  TC_Constant # (.UUID(64'd2159418541358820159 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_6 (.out(wire_4));
  TC_Constant # (.UUID(64'd3865030967482760074 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100)) Constant64_7 (.out(wire_65));
  TC_Shl # (.UUID(64'd256840837460643515 ^ UUID), .BIT_WIDTH(64'd64)) Shl64_8 (.in(wire_65), .shift(wire_63), .out(wire_25));
  TC_Add # (.UUID(64'd2069450991047535688 ^ UUID), .BIT_WIDTH(64'd8)) Add8_9 (.in0(wire_88), .in1(wire_48), .ci(1'd0), .out(wire_63), .co());
  TC_Constant # (.UUID(64'd890068480924790415 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_10 (.out(wire_1));
  TC_Mul # (.UUID(64'd1392401372469684178 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_11 (.in0(wire_51), .in1(wire_1), .out0(wire_88), .out1());
  TC_Constant # (.UUID(64'd2849228403424780629 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h8)) Constant32_12 (.out(wire_24));
  TC_Or # (.UUID(64'd2449338929424116540 ^ UUID), .BIT_WIDTH(64'd64)) Or64_13 (.in0(wire_72), .in1(wire_36), .out(wire_54));
  TC_Constant # (.UUID(64'd1543423362108290125 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h100000000000000)) Constant64_14 (.out(wire_74));
  TC_Equal # (.UUID(64'd4163658842919617091 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_15 (.in0(wire_9), .in1(wire_96), .out(wire_99));
  TC_Constant # (.UUID(64'd2675462162887539169 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h1800)) Constant32_16 (.out(wire_96));
  TC_Mux # (.UUID(64'd1930168901414496793 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_17 (.sel(wire_3), .in0(wire_100), .in1(wire_21[7:0]), .out(wire_80));
  TC_Switch # (.UUID(64'd2050260038134492089 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_18 (.en(wire_97), .in(wire_25), .out(wire_72));
  TC_Switch # (.UUID(64'd4459812316626182275 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_37), .in(wire_0), .out(wire_81));
  TC_Maker8 # (.UUID(64'd3476275697879983087 ^ UUID)) Maker8_20 (.in0(wire_17), .in1(wire_98), .in2(wire_91), .in3(wire_86), .in4(wire_53), .in5(wire_7), .in6(wire_39), .in7(wire_56), .out(wire_100));
  TC_Splitter8 # (.UUID(64'd2521255541794198669 ^ UUID)) Splitter8_21 (.in(wire_80), .out0(wire_37), .out1(wire_92), .out2(wire_55), .out3(wire_94), .out4(wire_46), .out5(wire_82), .out6(wire_50), .out7(wire_85));
  TC_Switch # (.UUID(64'd3245081307199932182 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_92), .in(wire_0), .out(wire_52));
  TC_Switch # (.UUID(64'd2002688052549140963 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_23 (.en(wire_55), .in(wire_0), .out(wire_49));
  TC_Switch # (.UUID(64'd107481461216313517 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_24 (.en(wire_94), .in(wire_0), .out(wire_15));
  TC_Splitter8 # (.UUID(64'd4255826572476153746 ^ UUID)) Splitter8_25 (.in(wire_59), .out0(wire_69), .out1(wire_45), .out2(wire_67), .out3(wire_11), .out4(wire_78), .out5(wire_95), .out6(wire_29), .out7(wire_84));
  TC_Switch # (.UUID(64'd1461177450814591256 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_26 (.en(wire_69), .in(wire_8), .out(wire_57));
  TC_Switch # (.UUID(64'd695816634534987300 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_27 (.en(wire_45), .in(wire_8), .out(wire_30));
  TC_Switch # (.UUID(64'd605369638144148965 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_28 (.en(wire_67), .in(wire_8), .out(wire_32));
  TC_Switch # (.UUID(64'd2158440079378329418 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_29 (.en(wire_11), .in(wire_8), .out(wire_33));
  TC_Switch # (.UUID(64'd1822975782747076870 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_30 (.en(wire_78), .in(wire_8), .out(wire_19));
  TC_Switch # (.UUID(64'd3972289372125110072 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_31 (.en(wire_95), .in(wire_8), .out(wire_18));
  TC_Switch # (.UUID(64'd4087363548528799060 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_32 (.en(wire_29), .in(wire_8), .out(wire_27));
  TC_Switch # (.UUID(64'd4071004930069955186 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_33 (.en(wire_84), .in(wire_8), .out(wire_61));
  TC_Not # (.UUID(64'd2063551563544788031 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_3), .out(wire_97));
  TC_Constant # (.UUID(64'd1477301682282254823 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h1)) Constant32_35 (.out(wire_89));
  TC_Or # (.UUID(64'd2383100013357812160 ^ UUID), .BIT_WIDTH(64'd32)) Or32_36 (.in0(wire_76), .in1(wire_89), .out(wire_8));
  TC_Shl # (.UUID(64'd1931844054005619464 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_37 (.in(wire_70), .shift(wire_24[7:0]), .out(wire_76));
  TC_Constant # (.UUID(64'd1647720820541862327 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h1)) Constant32_38 (.out(wire_68));
  TC_Or # (.UUID(64'd4577658088330867745 ^ UUID), .BIT_WIDTH(64'd64)) Or64_39 (.in0(wire_54), .in1({{32{1'b0}}, wire_68 }), .out(wire_0));
  TC_Switch # (.UUID(64'd1105450258378979929 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_40 (.en(wire_3), .in(wire_74), .out(wire_36));
  TC_Switch # (.UUID(64'd3633178823871315022 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_75), .in(wire_99), .out(wire_3));
  TC_Switch # (.UUID(64'd2715234750164652225 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_42 (.en(wire_46), .in(wire_0), .out(wire_34));
  TC_Switch # (.UUID(64'd1703957103141682707 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_43 (.en(wire_82), .in(wire_0), .out(wire_41));
  TC_Switch # (.UUID(64'd3116247898275579677 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_44 (.en(wire_50), .in(wire_0), .out(wire_13));
  TC_Switch # (.UUID(64'd1886574100080780526 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_45 (.en(wire_85), .in(wire_0), .out(wire_28));
  TC_Constant # (.UUID(64'd1716300220336083549 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hFFFF)) Constant16_46 (.out(wire_21));
  TC_Mux # (.UUID(64'd2070625018299700787 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_47 (.sel(wire_3), .in0(wire_66), .in1(wire_21), .out(wire_20));
  TC_Not # (.UUID(64'd4098144234192782196 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_22), .out(wire_90));
  TC_Constant # (.UUID(64'd3385451059797225464 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_49 (.out(wire_2));
  TC_Shl # (.UUID(64'd4330698639726977865 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_50 (.in(wire_2), .shift(wire_35), .out(wire_73));
  TC_Switch # (.UUID(64'd484212059188064426 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_51 (.en(wire_90), .in(wire_73), .out(wire_66));
  TC_Splitter8 # (.UUID(64'd335990418435108769 ^ UUID)) Splitter8_52 (.in(wire_64), .out0(wire_79), .out1(wire_38), .out2(wire_5), .out3(wire_62), .out4(wire_71), .out5(wire_6), .out6(wire_87), .out7(wire_93));
  TC_Switch # (.UUID(64'd1686490303216320774 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_53 (.en(wire_79), .in(wire_8), .out(wire_83));
  TC_Switch # (.UUID(64'd3394474682486717869 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_54 (.en(wire_38), .in(wire_8), .out(wire_40));
  TC_Switch # (.UUID(64'd3453098892598527541 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_55 (.en(wire_5), .in(wire_8), .out(wire_47));
  TC_Switch # (.UUID(64'd1969313976998410780 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_56 (.en(wire_62), .in(wire_8), .out(wire_16));
  TC_Switch # (.UUID(64'd736854851732662637 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_57 (.en(wire_71), .in(wire_8), .out(wire_26));
  TC_Switch # (.UUID(64'd305341364590474780 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_58 (.en(wire_6), .in(wire_8), .out(wire_14));
  TC_Switch # (.UUID(64'd3274241556523413121 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_59 (.en(wire_87), .in(wire_8), .out(wire_58));
  TC_Switch # (.UUID(64'd2925559771953586588 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_60 (.en(wire_93), .in(wire_8), .out(wire_44));
  TC_Splitter16 # (.UUID(64'd703182031863533036 ^ UUID)) Splitter16_61 (.in(wire_20), .out0(wire_59), .out1(wire_64));
  TC_Mul # (.UUID(64'd3291077814889728828 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_62 (.in0(wire_60[7:0]), .in1(wire_10), .out0(wire_31), .out1(wire_51));
  TC_Mul # (.UUID(64'd3820707656544130399 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_63 (.in0(wire_43[7:0]), .in1(wire_4), .out0(wire_35), .out1(wire_48));

  wire [63:0] wire_0;
  wire [7:0] wire_1;
  wire [15:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [31:0] wire_8;
  wire [31:0] wire_9;
  assign wire_9 = Address;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [63:0] wire_13;
  assign Output_23 = wire_13;
  wire [31:0] wire_14;
  assign Output_14 = wire_14;
  wire [63:0] wire_15;
  assign Output_20 = wire_15;
  wire [31:0] wire_16;
  assign Output_12 = wire_16;
  wire [0:0] wire_17;
  wire [31:0] wire_18;
  assign Output_6 = wire_18;
  wire [31:0] wire_19;
  assign Output_5 = wire_19;
  wire [15:0] wire_20;
  wire [15:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [31:0] wire_24;
  wire [63:0] wire_25;
  wire [31:0] wire_26;
  assign Output_13 = wire_26;
  wire [31:0] wire_27;
  assign Output_7 = wire_27;
  wire [63:0] wire_28;
  assign Output_24 = wire_28;
  wire [0:0] wire_29;
  wire [31:0] wire_30;
  assign Output_2 = wire_30;
  wire [7:0] wire_31;
  wire [31:0] wire_32;
  assign Output_3 = wire_32;
  wire [31:0] wire_33;
  assign Output_4 = wire_33;
  wire [63:0] wire_34;
  assign Output_21 = wire_34;
  wire [7:0] wire_35;
  wire [63:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [31:0] wire_40;
  assign Output_10 = wire_40;
  wire [63:0] wire_41;
  assign Output_22 = wire_41;
  wire [0:0] wire_42;
  wire [31:0] wire_43;
  wire [31:0] wire_44;
  assign Output_16 = wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [31:0] wire_47;
  assign Output_11 = wire_47;
  wire [7:0] wire_48;
  wire [63:0] wire_49;
  assign Output_19 = wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [63:0] wire_52;
  assign Output_18 = wire_52;
  wire [0:0] wire_53;
  wire [63:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [31:0] wire_57;
  assign Output_1 = wire_57;
  wire [31:0] wire_58;
  assign Output_15 = wire_58;
  wire [7:0] wire_59;
  wire [31:0] wire_60;
  wire [31:0] wire_61;
  assign Output_8 = wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [7:0] wire_64;
  wire [63:0] wire_65;
  wire [15:0] wire_66;
  wire [0:0] wire_67;
  wire [31:0] wire_68;
  wire [0:0] wire_69;
  wire [31:0] wire_70;
  assign wire_70 = Value;
  wire [0:0] wire_71;
  wire [63:0] wire_72;
  wire [15:0] wire_73;
  wire [63:0] wire_74;
  wire [0:0] wire_75;
  assign wire_75 = Enable;
  wire [31:0] wire_76;
  wire [31:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [7:0] wire_80;
  wire [63:0] wire_81;
  assign Output_17 = wire_81;
  wire [0:0] wire_82;
  wire [31:0] wire_83;
  assign Output_9 = wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [7:0] wire_88;
  wire [31:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [31:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [7:0] wire_100;

endmodule
