module _4bit_Decoder (clk, rst, \1_1 , \2_1 , \4_1 , \8_1 , \7 , \11 , \3 , \15 , \6 , \8_2 , \5 , \9 , \10 , \4_2 , \12 , \13 , \14 , \2_2 , \1_2 , \0 );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] \1_1 ;
  input  wire [0:0] \2_1 ;
  input  wire [0:0] \4_1 ;
  input  wire [0:0] \8_1 ;
  output  wire [0:0] \7 ;
  output  wire [0:0] \11 ;
  output  wire [0:0] \3 ;
  output  wire [0:0] \15 ;
  output  wire [0:0] \6 ;
  output  wire [0:0] \8_2 ;
  output  wire [0:0] \5 ;
  output  wire [0:0] \9 ;
  output  wire [0:0] \10 ;
  output  wire [0:0] \4_2 ;
  output  wire [0:0] \12 ;
  output  wire [0:0] \13 ;
  output  wire [0:0] \14 ;
  output  wire [0:0] \2_2 ;
  output  wire [0:0] \1_2 ;
  output  wire [0:0] \0 ;

  TC_And3 # (.UUID(64'd631691880289895914 ^ UUID), .BIT_WIDTH(64'd1)) And3_0 (.in0(wire_60), .in1(wire_16), .in2(wire_56), .out(wire_32));
  TC_And # (.UUID(64'd570263192918881500 ^ UUID), .BIT_WIDTH(64'd1)) And_1 (.in0(wire_53), .in1(wire_50), .out(wire_60));
  TC_Not # (.UUID(64'd4055959480987982074 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_7), .out(wire_53));
  TC_Not # (.UUID(64'd504647261216695913 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_2), .out(wire_50));
  TC_Not # (.UUID(64'd4464546700307020499 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_6), .out(wire_16));
  TC_Not # (.UUID(64'd87826712391748840 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_4), .out(wire_56));
  TC_And3 # (.UUID(64'd3437650392345874692 ^ UUID), .BIT_WIDTH(64'd1)) And3_6 (.in0(wire_80), .in1(wire_13), .in2(wire_46), .out(wire_74));
  TC_And # (.UUID(64'd2734826135142314724 ^ UUID), .BIT_WIDTH(64'd1)) And_7 (.in0(wire_7), .in1(wire_65), .out(wire_80));
  TC_Not # (.UUID(64'd3636390598591512326 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_6), .out(wire_13));
  TC_Not # (.UUID(64'd772683298208068349 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_4), .out(wire_46));
  TC_Not # (.UUID(64'd3720093155665021630 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_2), .out(wire_65));
  TC_And3 # (.UUID(64'd3468100056999563378 ^ UUID), .BIT_WIDTH(64'd1)) And3_11 (.in0(wire_57), .in1(wire_69), .in2(wire_41), .out(wire_19));
  TC_And # (.UUID(64'd1846765807919374199 ^ UUID), .BIT_WIDTH(64'd1)) And_12 (.in0(wire_54), .in1(wire_2), .out(wire_57));
  TC_Not # (.UUID(64'd3944775958458564079 ^ UUID), .BIT_WIDTH(64'd1)) Not_13 (.in(wire_7), .out(wire_54));
  TC_Not # (.UUID(64'd1355787431147599723 ^ UUID), .BIT_WIDTH(64'd1)) Not_14 (.in(wire_6), .out(wire_69));
  TC_Not # (.UUID(64'd2455930481895824666 ^ UUID), .BIT_WIDTH(64'd1)) Not_15 (.in(wire_4), .out(wire_41));
  TC_And3 # (.UUID(64'd2920462676885562663 ^ UUID), .BIT_WIDTH(64'd1)) And3_16 (.in0(wire_52), .in1(wire_48), .in2(wire_85), .out(wire_99));
  TC_And # (.UUID(64'd4167424231857602842 ^ UUID), .BIT_WIDTH(64'd1)) And_17 (.in0(wire_7), .in1(wire_2), .out(wire_52));
  TC_Not # (.UUID(64'd1756443747051396474 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_6), .out(wire_48));
  TC_Not # (.UUID(64'd3318056850283048249 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_4), .out(wire_85));
  TC_And3 # (.UUID(64'd2569057375939886449 ^ UUID), .BIT_WIDTH(64'd1)) And3_20 (.in0(wire_90), .in1(wire_6), .in2(wire_21), .out(wire_26));
  TC_And # (.UUID(64'd1968058018053543343 ^ UUID), .BIT_WIDTH(64'd1)) And_21 (.in0(wire_20), .in1(wire_15), .out(wire_90));
  TC_Not # (.UUID(64'd4149321274639640752 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_7), .out(wire_20));
  TC_Not # (.UUID(64'd1566567313842736592 ^ UUID), .BIT_WIDTH(64'd1)) Not_23 (.in(wire_2), .out(wire_15));
  TC_Not # (.UUID(64'd1836063106694412281 ^ UUID), .BIT_WIDTH(64'd1)) Not_24 (.in(wire_4), .out(wire_21));
  TC_And3 # (.UUID(64'd4334170431590759070 ^ UUID), .BIT_WIDTH(64'd1)) And3_25 (.in0(wire_61), .in1(wire_6), .in2(wire_36), .out(wire_95));
  TC_And # (.UUID(64'd415083169861684526 ^ UUID), .BIT_WIDTH(64'd1)) And_26 (.in0(wire_7), .in1(wire_5), .out(wire_61));
  TC_Not # (.UUID(64'd1134923669678933276 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_2), .out(wire_5));
  TC_Not # (.UUID(64'd2886678207462735138 ^ UUID), .BIT_WIDTH(64'd1)) Not_28 (.in(wire_4), .out(wire_36));
  TC_And3 # (.UUID(64'd188062065042578749 ^ UUID), .BIT_WIDTH(64'd1)) And3_29 (.in0(wire_76), .in1(wire_6), .in2(wire_66), .out(wire_45));
  TC_And # (.UUID(64'd2460638328327494292 ^ UUID), .BIT_WIDTH(64'd1)) And_30 (.in0(wire_71), .in1(wire_2), .out(wire_76));
  TC_Not # (.UUID(64'd3900559227156551805 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_7), .out(wire_71));
  TC_Not # (.UUID(64'd2997939628519448689 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_4), .out(wire_66));
  TC_And3 # (.UUID(64'd974378858837864169 ^ UUID), .BIT_WIDTH(64'd1)) And3_33 (.in0(wire_91), .in1(wire_6), .in2(wire_28), .out(wire_11));
  TC_And # (.UUID(64'd425178247384331206 ^ UUID), .BIT_WIDTH(64'd1)) And_34 (.in0(wire_7), .in1(wire_2), .out(wire_91));
  TC_Not # (.UUID(64'd4380552074478123722 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_4), .out(wire_28));
  TC_And3 # (.UUID(64'd896788497510746464 ^ UUID), .BIT_WIDTH(64'd1)) And3_36 (.in0(wire_79), .in1(wire_38), .in2(wire_4), .out(wire_73));
  TC_And # (.UUID(64'd3938047067186107761 ^ UUID), .BIT_WIDTH(64'd1)) And_37 (.in0(wire_37), .in1(wire_77), .out(wire_79));
  TC_Not # (.UUID(64'd73163863177738551 ^ UUID), .BIT_WIDTH(64'd1)) Not_38 (.in(wire_7), .out(wire_37));
  TC_Not # (.UUID(64'd3380687016328036699 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_2), .out(wire_77));
  TC_Not # (.UUID(64'd1365874160878312651 ^ UUID), .BIT_WIDTH(64'd1)) Not_40 (.in(wire_6), .out(wire_38));
  TC_And3 # (.UUID(64'd1897297487657023211 ^ UUID), .BIT_WIDTH(64'd1)) And3_41 (.in0(wire_49), .in1(wire_62), .in2(wire_4), .out(wire_63));
  TC_And # (.UUID(64'd1258527878262494242 ^ UUID), .BIT_WIDTH(64'd1)) And_42 (.in0(wire_7), .in1(wire_9), .out(wire_49));
  TC_Not # (.UUID(64'd3464705032636047656 ^ UUID), .BIT_WIDTH(64'd1)) Not_43 (.in(wire_2), .out(wire_9));
  TC_Not # (.UUID(64'd3473152955628639238 ^ UUID), .BIT_WIDTH(64'd1)) Not_44 (.in(wire_6), .out(wire_62));
  TC_And3 # (.UUID(64'd2783289211952775351 ^ UUID), .BIT_WIDTH(64'd1)) And3_45 (.in0(wire_92), .in1(wire_98), .in2(wire_4), .out(wire_64));
  TC_And # (.UUID(64'd2347315004226464140 ^ UUID), .BIT_WIDTH(64'd1)) And_46 (.in0(wire_10), .in1(wire_2), .out(wire_92));
  TC_Not # (.UUID(64'd2893048661734952089 ^ UUID), .BIT_WIDTH(64'd1)) Not_47 (.in(wire_7), .out(wire_10));
  TC_Not # (.UUID(64'd2027922108154434464 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_6), .out(wire_98));
  TC_And3 # (.UUID(64'd2210692075283983171 ^ UUID), .BIT_WIDTH(64'd1)) And3_49 (.in0(wire_14), .in1(wire_72), .in2(wire_4), .out(wire_75));
  TC_And # (.UUID(64'd750893363983607753 ^ UUID), .BIT_WIDTH(64'd1)) And_50 (.in0(wire_7), .in1(wire_2), .out(wire_14));
  TC_Not # (.UUID(64'd1308304970739126268 ^ UUID), .BIT_WIDTH(64'd1)) Not_51 (.in(wire_6), .out(wire_72));
  TC_And3 # (.UUID(64'd2077791055199310333 ^ UUID), .BIT_WIDTH(64'd1)) And3_52 (.in0(wire_59), .in1(wire_6), .in2(wire_4), .out(wire_58));
  TC_And # (.UUID(64'd3396760489957176935 ^ UUID), .BIT_WIDTH(64'd1)) And_53 (.in0(wire_27), .in1(wire_94), .out(wire_59));
  TC_Not # (.UUID(64'd3497892084035099871 ^ UUID), .BIT_WIDTH(64'd1)) Not_54 (.in(wire_7), .out(wire_27));
  TC_Not # (.UUID(64'd4322149666828256789 ^ UUID), .BIT_WIDTH(64'd1)) Not_55 (.in(wire_2), .out(wire_94));
  TC_And3 # (.UUID(64'd4130284332433004246 ^ UUID), .BIT_WIDTH(64'd1)) And3_56 (.in0(wire_83), .in1(wire_6), .in2(wire_4), .out(wire_29));
  TC_And # (.UUID(64'd242325210640456277 ^ UUID), .BIT_WIDTH(64'd1)) And_57 (.in0(wire_7), .in1(wire_25), .out(wire_83));
  TC_Not # (.UUID(64'd1551208013100794203 ^ UUID), .BIT_WIDTH(64'd1)) Not_58 (.in(wire_2), .out(wire_25));
  TC_And3 # (.UUID(64'd786451316106540696 ^ UUID), .BIT_WIDTH(64'd1)) And3_59 (.in0(wire_93), .in1(wire_6), .in2(wire_4), .out(wire_0));
  TC_And # (.UUID(64'd191331196645785238 ^ UUID), .BIT_WIDTH(64'd1)) And_60 (.in0(wire_39), .in1(wire_2), .out(wire_93));
  TC_Not # (.UUID(64'd2013225323766124818 ^ UUID), .BIT_WIDTH(64'd1)) Not_61 (.in(wire_7), .out(wire_39));
  TC_And3 # (.UUID(64'd4421779969158748059 ^ UUID), .BIT_WIDTH(64'd1)) And3_62 (.in0(wire_82), .in1(wire_6), .in2(wire_4), .out(wire_88));
  TC_And # (.UUID(64'd1785139406016315052 ^ UUID), .BIT_WIDTH(64'd1)) And_63 (.in0(wire_7), .in1(wire_2), .out(wire_82));
  TC_Switch # (.UUID(64'd3034604376454019258 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_64 (.en(wire_32), .in(wire_70), .out(wire_8));
  TC_Constant # (.UUID(64'd1288316162819049283 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_65 (.out(wire_70));
  TC_Switch # (.UUID(64'd790256782469417320 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_74), .in(wire_18), .out(wire_67));
  TC_Constant # (.UUID(64'd1611432490062290311 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_67 (.out(wire_18));
  TC_Switch # (.UUID(64'd4418756422035915438 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_68 (.en(wire_19), .in(wire_43), .out(wire_68));
  TC_Constant # (.UUID(64'd336023926348934563 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_69 (.out(wire_43));
  TC_Switch # (.UUID(64'd1415791970800101993 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_70 (.en(wire_99), .in(wire_1), .out(wire_3));
  TC_Constant # (.UUID(64'd3000239064114474112 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_71 (.out(wire_1));
  TC_Switch # (.UUID(64'd3511636667321256480 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_72 (.en(wire_26), .in(wire_34), .out(wire_51));
  TC_Constant # (.UUID(64'd675924624058025154 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_73 (.out(wire_34));
  TC_Switch # (.UUID(64'd3901122780939301375 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_74 (.en(wire_95), .in(wire_42), .out(wire_40));
  TC_Constant # (.UUID(64'd4164162661660036947 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_75 (.out(wire_42));
  TC_Switch # (.UUID(64'd1635843679600751182 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_76 (.en(wire_45), .in(wire_33), .out(wire_30));
  TC_Constant # (.UUID(64'd3343297195376566013 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_77 (.out(wire_33));
  TC_Switch # (.UUID(64'd120029340335375031 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_78 (.en(wire_11), .in(wire_22), .out(wire_44));
  TC_Constant # (.UUID(64'd3699079282922615612 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_79 (.out(wire_22));
  TC_Switch # (.UUID(64'd2969442901624594062 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_80 (.en(wire_73), .in(wire_55), .out(wire_97));
  TC_Constant # (.UUID(64'd3524771667935717177 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_81 (.out(wire_55));
  TC_Switch # (.UUID(64'd770322839737333588 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_82 (.en(wire_63), .in(wire_84), .out(wire_89));
  TC_Constant # (.UUID(64'd1472050705962282008 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_83 (.out(wire_84));
  TC_Switch # (.UUID(64'd783698755752463085 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_84 (.en(wire_64), .in(wire_35), .out(wire_78));
  TC_Constant # (.UUID(64'd360966707612435960 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_85 (.out(wire_35));
  TC_Switch # (.UUID(64'd3908323290067766716 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_86 (.en(wire_75), .in(wire_87), .out(wire_24));
  TC_Constant # (.UUID(64'd2693169534973350234 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_87 (.out(wire_87));
  TC_Switch # (.UUID(64'd4147170937949799501 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_88 (.en(wire_58), .in(wire_47), .out(wire_31));
  TC_Constant # (.UUID(64'd1968099585390582827 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_89 (.out(wire_47));
  TC_Switch # (.UUID(64'd3625912546760542287 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_90 (.en(wire_29), .in(wire_23), .out(wire_96));
  TC_Constant # (.UUID(64'd1357270235827237278 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_91 (.out(wire_23));
  TC_Switch # (.UUID(64'd3134605850462075464 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_92 (.en(wire_0), .in(wire_81), .out(wire_17));
  TC_Constant # (.UUID(64'd3086641151123060984 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_93 (.out(wire_81));
  TC_Switch # (.UUID(64'd3457539279353942043 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_94 (.en(wire_88), .in(wire_12), .out(wire_86));
  TC_Constant # (.UUID(64'd354868037566896794 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_95 (.out(wire_12));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign wire_2 = \2_1 ;
  wire [0:0] wire_3;
  assign \3  = wire_3;
  wire [0:0] wire_4;
  assign wire_4 = \8_1 ;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  assign wire_6 = \4_1 ;
  wire [0:0] wire_7;
  assign wire_7 = \1_1 ;
  wire [0:0] wire_8;
  assign \0  = wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  assign \14  = wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  assign \11  = wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  assign \6  = wire_30;
  wire [0:0] wire_31;
  assign \12  = wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  assign \5  = wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  assign \7  = wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  assign \4_2  = wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  assign \1_2  = wire_67;
  wire [0:0] wire_68;
  assign \2_2  = wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  assign \10  = wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  assign \15  = wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  assign \9  = wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  assign \13  = wire_96;
  wire [0:0] wire_97;
  assign \8_2  = wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;

endmodule
