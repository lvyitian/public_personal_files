module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_1), .en(wire_75), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_34), .in(arch_input_value), .out(wire_20));
  TC_Program8_4 # (.UUID(64'd4489305393227859486 ^ UUID), .DEFAULT_FILE_NAME("Program8_4_3E4D37784397861E.w8.bin"), .ARG_SIG("Program8_4_3E4D37784397861E=%s")) Program8_4_2 (.clk(clk), .rst(rst), .address(wire_53), .out0(wire_22), .out1(wire_65), .out2(wire_54), .out3(wire_73));
  TC_Counter # (.UUID(64'd1175999672554394000 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_3 (.clk(clk), .rst(rst), .save(wire_9), .in(wire_1), .out(wire_53));
  TC_Splitter8 # (.UUID(64'd3496280010280654809 ^ UUID)) Splitter8_4 (.in(wire_92), .out0(wire_21), .out1(wire_30), .out2(wire_23), .out3(wire_88), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1350359362790102949 ^ UUID)) Splitter8_5 (.in(wire_19), .out0(wire_61), .out1(wire_83), .out2(wire_81), .out3(wire_59), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3688384451292696869 ^ UUID)) Splitter8_6 (.in(wire_52), .out0(wire_76), .out1(wire_6), .out2(wire_69), .out3(wire_35), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3357720912797461292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_55), .in(wire_53), .out());
  TC_Maker8 # (.UUID(64'd2922775923237819214 ^ UUID)) Maker8_8 (.in0(wire_90), .in1(wire_63), .in2(wire_32), .in3(wire_58), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_74));
  TC_Splitter8 # (.UUID(64'd4136660363423911410 ^ UUID)) Splitter8_9 (.in(wire_22), .out0(wire_90), .out1(wire_63), .out2(wire_32), .out3(wire_58), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd4550958897663313502 ^ UUID)) Splitter8_10 (.in(wire_22), .out0(wire_51), .out1(wire_64), .out2(wire_29), .out3(wire_71), .out4(wire_93), .out5(wire_26), .out6(wire_46), .out7(wire_68));
  TC_Maker8 # (.UUID(64'd3153840370766490713 ^ UUID)) Maker8_11 (.in0(wire_51), .in1(wire_64), .in2(wire_29), .in3(wire_71), .in4(wire_93), .in5(wire_26), .in6(wire_46), .in7(wire_68), .out(wire_37));
  TC_Constant # (.UUID(64'd4029987529778329422 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out(wire_82));
  TC_Constant # (.UUID(64'd47372170638122597 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_11));
  TC_Constant # (.UUID(64'd3010400910295959985 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_89));
  TC_Constant # (.UUID(64'd1353887318054096472 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out(wire_25));
  TC_Constant # (.UUID(64'd4461919415197064488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_44));
  TC_Constant # (.UUID(64'd2551986311311524963 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out(wire_45));
  TC_Switch # (.UUID(64'd201407107924193690 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_87), .in(wire_42), .out(wire_10_5));
  TC_Switch # (.UUID(64'd3784926049681585699 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_95), .in(wire_42), .out(wire_8_5));
  TC_Switch # (.UUID(64'd3418942253385023549 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_94), .in(wire_27), .out(wire_10_1));
  TC_Switch # (.UUID(64'd3104771108315787100 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_85), .in(wire_27), .out(wire_8_6));
  TC_Switch # (.UUID(64'd494263610589549334 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_47), .in(wire_0), .out(wire_10_3));
  TC_Switch # (.UUID(64'd4455028313033582898 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_39), .in(wire_0), .out(wire_8_4));
  TC_Switch # (.UUID(64'd977062972681925203 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_49), .in(wire_4), .out(wire_10_4));
  TC_Switch # (.UUID(64'd2935373336597064260 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_14), .in(wire_4), .out(wire_8_0));
  TC_Switch # (.UUID(64'd2595310988575568445 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_28), .in(wire_48), .out(wire_10_2));
  TC_Switch # (.UUID(64'd3649926646471230167 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_50), .in(wire_48), .out(wire_8_3));
  TC_Switch # (.UUID(64'd115863760055946247 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_67), .in(wire_62), .out(wire_10_0));
  TC_Switch # (.UUID(64'd459043271910661458 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_91), .in(wire_62), .out(wire_8_1));
  TC_Switch # (.UUID(64'd4275937720180353902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_40), .in(wire_53), .out());
  TC_Switch # (.UUID(64'd2718446434835356700 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_38), .in(wire_20), .out(wire_10_6));
  TC_Switch # (.UUID(64'd1811299859375739998 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_79), .in(wire_20), .out(wire_8_2));
  TC_Or # (.UUID(64'd117421755651659184 ^ UUID), .BIT_WIDTH(64'd1)) Or_33 (.in0(wire_38), .in1(wire_79), .out(wire_34));
  TC_Switch # (.UUID(64'd262409980643160938 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_31), .in(wire_54), .out(wire_8_9));
  TC_Switch # (.UUID(64'd2764614579549035605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_60), .in(wire_65), .out(wire_10_8));
  TC_Switch # (.UUID(64'd2974460371787013801 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_24), .in(wire_41), .out(wire_1_0));
  TC_Mux # (.UUID(64'd1769789085559769130 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_37 (.sel(wire_31), .in0(wire_54), .in1(wire_15), .out(wire_19));
  TC_Mux # (.UUID(64'd1404337327044278632 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_60), .in0(wire_65), .in1(wire_13), .out(wire_92));
  TC_Constant # (.UUID(64'd4387708643330744374 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_39 (.out(wire_13));
  TC_Constant # (.UUID(64'd2430039925245603401 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_40 (.out(wire_15));
  TC_Switch # (.UUID(64'd3877536405880520929 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_72), .in(wire_80), .out(wire_16));
  TC_Constant # (.UUID(64'd2430392602802046886 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_42 (.out(wire_84));
  TC_Mux # (.UUID(64'd1559488034901936773 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_43 (.sel(wire_16), .in0(wire_73), .in1(wire_84), .out(wire_52));
  TC_Switch # (.UUID(64'd3981948550050450551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_16), .in(wire_73), .out(wire_1_1));
  TC_Ram # (.UUID(64'd1683242105781375453 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_45 (.clk(clk), .rst(rst), .load(wire_77), .save(wire_78), .address({{24{1'b0}}, wire_18 }), .in0({{56{1'b0}}, wire_1 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_57), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd1949247607308932292 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_46 (.out(wire_5));
  TC_Or # (.UUID(64'd2571069615494455195 ^ UUID), .BIT_WIDTH(64'd1)) Or_47 (.in0(wire_33), .in1(wire_43), .out(wire_77));
  TC_Switch # (.UUID(64'd3896516251333244950 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_56), .in(wire_70), .out(wire_10_7));
  TC_Switch # (.UUID(64'd4219278115069450234 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_86), .in(wire_70), .out(wire_8_7));
  TC_Switch # (.UUID(64'd875265095609107539 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_33), .in(wire_57[7:0]), .out(wire_10_9));
  TC_Switch # (.UUID(64'd1025433274855748469 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_43), .in(wire_57[7:0]), .out(wire_8_8));
  _4bit_Decoder # (.UUID(64'd188593635878702660 ^ UUID)) _4bit_Decoder_52 (.clk(clk), .rst(rst), .\1_1 (wire_21), .\2_1 (wire_30), .\4_1 (wire_23), .\8_1 (wire_88), .\7 (wire_38), .\11 (), .\3 (wire_49), .\15 (), .\6 (wire_55), .\8_2 (wire_56), .\5 (wire_67), .\9 (wire_33), .\10 (), .\4_2 (wire_28), .\12 (), .\13 (), .\14 (), .\2_2 (wire_47), .\1_2 (wire_94), .\0 (wire_87));
  _4bit_Decoder # (.UUID(64'd3657203059375966986 ^ UUID)) _4bit_Decoder_53 (.clk(clk), .rst(rst), .\1_1 (wire_61), .\2_1 (wire_83), .\4_1 (wire_81), .\8_1 (wire_59), .\7 (wire_79), .\11 (), .\3 (wire_14), .\15 (), .\6 (wire_40), .\8_2 (wire_86), .\5 (wire_91), .\9 (wire_43), .\10 (), .\4_2 (wire_50), .\12 (), .\13 (), .\14 (), .\2_2 (wire_39), .\1_2 (wire_85), .\0 (wire_95));
  _4bit_Decoder # (.UUID(64'd4526675728054865805 ^ UUID)) _4bit_Decoder_54 (.clk(clk), .rst(rst), .\1_1 (wire_76), .\2_1 (wire_6), .\4_1 (wire_69), .\8_1 (wire_35), .\7 (wire_75), .\11 (), .\3 (wire_2), .\15 (), .\6 (wire_9), .\8_2 (wire_66), .\5 (wire_12), .\9 (wire_78), .\10 (), .\4_2 (wire_7), .\12 (), .\13 (), .\14 (), .\2_2 (wire_3), .\1_2 (wire_17), .\0 (wire_36));
  RegisterPlus # (.UUID(64'd1898575026262245003 ^ UUID)) RegisterPlus_55 (.clk(clk), .rst(rst), .\�_____ (wire_82), .\�___________ (wire_1), .\�_____ (wire_36), .\�___________ (), .Output(wire_42));
  RegisterPlus # (.UUID(64'd201486149512558618 ^ UUID)) RegisterPlus_56 (.clk(clk), .rst(rst), .\�_____ (wire_11), .\�___________ (wire_1), .\�_____ (wire_17), .\�___________ (), .Output(wire_27));
  RegisterPlus # (.UUID(64'd4130910523704063521 ^ UUID)) RegisterPlus_57 (.clk(clk), .rst(rst), .\�_____ (wire_89), .\�___________ (wire_1), .\�_____ (wire_3), .\�___________ (), .Output(wire_0));
  RegisterPlus # (.UUID(64'd579904311903668382 ^ UUID)) RegisterPlus_58 (.clk(clk), .rst(rst), .\�_____ (wire_25), .\�___________ (wire_1), .\�_____ (wire_2), .\�___________ (), .Output(wire_4));
  RegisterPlus # (.UUID(64'd2026589517635316452 ^ UUID)) RegisterPlus_59 (.clk(clk), .rst(rst), .\�_____ (wire_44), .\�___________ (wire_1), .\�_____ (wire_7), .\�___________ (), .Output(wire_48));
  RegisterPlus # (.UUID(64'd1622410096212380183 ^ UUID)) RegisterPlus_60 (.clk(clk), .rst(rst), .\�_____ (wire_45), .\�___________ (wire_1), .\�_____ (wire_12), .\�___________ (), .Output(wire_62));
  LEG_ALU # (.UUID(64'd740631443788402157 ^ UUID)) LEG_ALU_61 (.clk(clk), .rst(rst), .\�_____ (wire_74), .\�______1 (wire_10), .\�______2 (wire_8), .Output(wire_41));
  LEG_COND # (.UUID(64'd999600516743479399 ^ UUID)) LEG_COND_62 (.clk(clk), .rst(rst), .ARG1(wire_10), .ARG2(wire_8), .\�_____ (wire_22), .Output(wire_80));
  RegisterPlus # (.UUID(64'd471658098348471390 ^ UUID)) RegisterPlus_63 (.clk(clk), .rst(rst), .\�_____ (wire_5), .\�___________ (wire_1), .\�_____ (wire_66), .\�___________ (wire_18), .Output(wire_70));
  LEG_DEC # (.UUID(64'd2015393024950033718 ^ UUID)) LEG_DEC_64 (.clk(clk), .rst(rst), .OPCODE(wire_37), .IMMEDIATE1(wire_60), .IMMEDIATE2(wire_31), .CALCULATION(wire_24), .JUMP(wire_72));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_8_0;
  wire [7:0] wire_8_1;
  wire [7:0] wire_8_2;
  wire [7:0] wire_8_3;
  wire [7:0] wire_8_4;
  wire [7:0] wire_8_5;
  wire [7:0] wire_8_6;
  wire [7:0] wire_8_7;
  wire [7:0] wire_8_8;
  wire [7:0] wire_8_9;
  assign wire_8 = wire_8_0|wire_8_1|wire_8_2|wire_8_3|wire_8_4|wire_8_5|wire_8_6|wire_8_7|wire_8_8|wire_8_9;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_10_0;
  wire [7:0] wire_10_1;
  wire [7:0] wire_10_2;
  wire [7:0] wire_10_3;
  wire [7:0] wire_10_4;
  wire [7:0] wire_10_5;
  wire [7:0] wire_10_6;
  wire [7:0] wire_10_7;
  wire [7:0] wire_10_8;
  wire [7:0] wire_10_9;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2|wire_10_3|wire_10_4|wire_10_5|wire_10_6|wire_10_7|wire_10_8|wire_10_9;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  assign arch_input_enable = wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [7:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [7:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [63:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [7:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [7:0] wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;
  assign arch_output_enable = wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [7:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;

endmodule
