module RISCzmV (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Ram # (.UUID(64'd98204067416641251 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd1030360)) Ram_0 (.clk(clk), .rst(rst), .load(wire_286), .save(wire_286), .address(wire_25[31:0]), .in0(wire_241), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_0), .out1(), .out2(), .out3());
  TC_FileLoader # (.UUID(64'd2878462717155625984 ^ UUID), .DEFAULT_FILE_NAME("turning-complete-riscv")) FileLoader_1 (.clk(clk), .rst(rst), .en(wire_133), .address(wire_414), .out(wire_323));
  TC_Register # (.UUID(64'd1203092348560168365 ^ UUID), .BIT_WIDTH(64'd64)) Register64_2 (.clk(clk), .rst(rst), .load(wire_165), .save(wire_153), .in(wire_323), .out(wire_66));
  TC_Equal # (.UUID(64'd3062847367553117909 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_3 (.in0(64'd0), .in1(wire_66), .out(wire_153));
  TC_Mux # (.UUID(64'd1930940828089793147 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_4 (.sel(wire_320), .in0(wire_136), .in1(wire_400), .out(wire_414));
  TC_Constant # (.UUID(64'd3380699531870645725 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_5 (.out(wire_136));
  TC_And # (.UUID(64'd1858582780564394731 ^ UUID), .BIT_WIDTH(64'd1)) And_6 (.in0(wire_210), .in1(wire_64), .out(wire_151));
  TC_Not # (.UUID(64'd1927697609643890799 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_153), .out(wire_210));
  TC_Constant # (.UUID(64'd4353625534986538219 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out(wire_165));
  TC_Not # (.UUID(64'd155787763123756012 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_153), .out(wire_320));
  TC_Not # (.UUID(64'd4583681398335491468 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_151), .out(wire_133));
  TC_Halt # (.UUID(64'd3915690226323091877 ^ UUID), .HALT_MESSAGE("Instruction Decoder Error")) Halt_11 (.clk(clk), .rst(rst), .en(wire_384));
  TC_Halt # (.UUID(64'd2599441231298045646 ^ UUID), .HALT_MESSAGE("ALU Error")) Halt_12 (.clk(clk), .rst(rst), .en(wire_395));
  TC_Or # (.UUID(64'd2434705228045369708 ^ UUID), .BIT_WIDTH(64'd1)) Or_13 (.in0(wire_317), .in1(wire_157), .out(wire_107));
  TC_Halt # (.UUID(64'd1082213053476870366 ^ UUID), .HALT_MESSAGE("Program Loaded")) Halt_14 (.clk(clk), .rst(rst), .en(1'd0));
  TC_DelayLine # (.UUID(64'd3290414157599741036 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_15 (.clk(clk), .rst(rst), .in(wire_151), .out(wire_349));
  TC_Xor # (.UUID(64'd3191129607970482768 ^ UUID), .BIT_WIDTH(64'd1)) Xor_16 (.in0(wire_349), .in1(wire_151), .out());
  TC_Constant # (.UUID(64'd310464359691240818 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h1000)) Constant32_17 (.out(wire_325));
  TC_Or # (.UUID(64'd3157666206962771571 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_153), .in1(wire_151), .out(wire_218));
  TC_Counter # (.UUID(64'd913859885921307876 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd8)) Counter64_19 (.clk(clk), .rst(rst), .save(wire_218), .in(wire_66), .out(wire_310));
  TC_Constant # (.UUID(64'd1803058630330213009 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h0)) Constant64_20 (.out(wire_232));
  TC_Add # (.UUID(64'd765698919337433620 ^ UUID), .BIT_WIDTH(64'd64)) Add64_21 (.in0(wire_310), .in1(wire_232), .ci(1'd0), .out(wire_400), .co());
  TC_LessU # (.UUID(64'd3522453922805080720 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_22 (.in0(wire_400), .in1(wire_66), .out(wire_226));
  TC_Not # (.UUID(64'd2083959471467750465 ^ UUID), .BIT_WIDTH(64'd1)) Not_23 (.in(wire_226), .out(wire_64));
  TC_And # (.UUID(64'd2384575025999119233 ^ UUID), .BIT_WIDTH(64'd1)) And_24 (.in0(wire_151), .in1(wire_182), .out(wire_373));
  TC_Mux # (.UUID(64'd4053199106919888041 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_25 (.sel(wire_356), .in0(wire_109[31:0]), .in1(wire_174), .out(wire_243));
  TC_Not # (.UUID(64'd2511006902236747738 ^ UUID), .BIT_WIDTH(64'd1)) Not_26 (.in(wire_182), .out(wire_356));
  TC_Or # (.UUID(64'd916758513425679763 ^ UUID), .BIT_WIDTH(64'd1)) Or_27 (.in0(wire_314), .in1(wire_90), .out(wire_317));
  TC_Mux # (.UUID(64'd2044231173657355104 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_28 (.sel(wire_151), .in0(wire_224), .in1(wire_108), .out(wire_231));
  TC_Mux # (.UUID(64'd2032211576538499296 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_29 (.sel(wire_151), .in0(wire_326), .in1(wire_306), .out(wire_115));
  TC_Constant # (.UUID(64'd686405128408528809 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_30 (.out(wire_224));
  TC_Constant # (.UUID(64'd2123028207882148082 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_31 (.out(wire_326));
  TC_Mux # (.UUID(64'd2721024215629092200 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_32 (.sel(wire_151), .in0(wire_310), .in1({{32{1'b0}}, wire_33 }), .out(wire_62));
  TC_Mux # (.UUID(64'd192770063111330505 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_33 (.sel(wire_151), .in0(wire_323), .in1({{32{1'b0}}, wire_1 }), .out(wire_9));
  TC_And # (.UUID(64'd3849349637502455647 ^ UUID), .BIT_WIDTH(64'd1)) And_34 (.in0(wire_151), .in1(wire_185), .out(wire_261));
  TC_Not # (.UUID(64'd993212363916678177 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_356), .out(wire_185));
  TC_Splitter32 # (.UUID(64'd1492107866582490488 ^ UUID)) Splitter32_36 (.in(wire_243), .out0(), .out1(), .out2(wire_217), .out3());
  TC_Splitter8 # (.UUID(64'd3327209537799980802 ^ UUID)) Splitter8_37 (.in(wire_217), .out0(), .out1(), .out2(), .out3(), .out4(wire_335), .out5(), .out6(), .out7());
  TC_Halt # (.UUID(64'd769548899855801389 ^ UUID), .HALT_MESSAGE("Test Failed")) Halt_38 (.clk(clk), .rst(rst), .en(wire_164));
  TC_And # (.UUID(64'd4286157878935432209 ^ UUID), .BIT_WIDTH(64'd1)) And_39 (.in0(wire_237), .in1(wire_335), .out(wire_164));
  TC_And # (.UUID(64'd3980779742889827357 ^ UUID), .BIT_WIDTH(64'd1)) And_40 (.in0(wire_237), .in1(wire_380), .out(wire_360));
  TC_Not # (.UUID(64'd977160974774792269 ^ UUID), .BIT_WIDTH(64'd1)) Not_41 (.in(wire_335), .out(wire_380));
  TC_Counter # (.UUID(64'd1389921540193080113 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_42 (.clk(clk), .rst(rst), .save(wire_391), .in(wire_329), .out(wire_329));
  TC_Not # (.UUID(64'd63554530343823950 ^ UUID), .BIT_WIDTH(64'd1)) Not_43 (.in(wire_360), .out(wire_391));
  TC_Console # (.UUID(64'd3687955947483314541 ^ UUID)) Console_44 (.clk(clk), .rst(rst), .offset(wire_293));
  TC_Constant # (.UUID(64'd3178684649331147699 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h400)) Constant32_45 (.out(wire_293));
  TC_Constant # (.UUID(64'd3399871130822417032 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h0)) Constant32_46 (.out(wire_448));
  TC_Equal # (.UUID(64'd550695988771256162 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_47 (.in0(wire_33), .in1(wire_448), .out(wire_440));
  TC_Halt # (.UUID(64'd2984768372604569257 ^ UUID), .HALT_MESSAGE("Breakpoint")) Halt_48 (.clk(clk), .rst(rst), .en(wire_440));
  TC_Switch # (.UUID(64'd1263814109437966602 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_49 (.en(wire_286), .in(wire_0), .out(wire_29_0));
  TC_LessU # (.UUID(64'd2726535354240853256 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_50 (.in0(wire_62), .in1(wire_345), .out(wire_286));
  TC_Constant # (.UUID(64'd1233951608221554714 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFF000000)) Constant64_51 (.out(wire_345));
  TC_Not # (.UUID(64'd1039692102739057368 ^ UUID), .BIT_WIDTH(64'd1)) Not_52 (.in(wire_286), .out(wire_36));
  TC_Equal # (.UUID(64'd1910671886081223482 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_53 (.in0(wire_62), .in1(wire_416), .out(wire_307));
  TC_Constant # (.UUID(64'd3670082939622378505 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFF000100)) Constant64_54 (.out(wire_416));
  TC_And # (.UUID(64'd3820054277743105768 ^ UUID), .BIT_WIDTH(64'd1)) And_55 (.in0(wire_36), .in1(wire_307), .out(wire_197));
  TC_Switch # (.UUID(64'd314070488467476831 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_56 (.en(wire_197), .in({{48{1'b0}}, wire_369 }), .out(wire_29_1));
  TC_Timing # (.UUID(64'd3367404360086462607 ^ UUID)) Timing_57 (.en(wire_370), .out(wire_29_2));
  TC_Equal # (.UUID(64'd396815649411487662 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_58 (.in0(wire_62), .in1(wire_98), .out(wire_212));
  TC_Constant # (.UUID(64'd632468375258568612 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFF000200)) Constant64_59 (.out(wire_98));
  TC_And # (.UUID(64'd3883096592534712930 ^ UUID), .BIT_WIDTH(64'd1)) And_60 (.in0(wire_36), .in1(wire_212), .out(wire_370));
  TC_Maker16 # (.UUID(64'd1967257727895694274 ^ UUID)) Maker16_61 (.in0({{7{1'b0}}, wire_268 }), .in1(wire_201), .out(wire_369));
  TC_Shl # (.UUID(64'd1589164205674529769 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_62 (.in({{7{1'b0}}, wire_337 }), .shift(wire_437), .out(wire_415));
  TC_Constant # (.UUID(64'd62967053956405745 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_63 (.out(wire_437));
  TC_Or # (.UUID(64'd416113240382239360 ^ UUID), .BIT_WIDTH(64'd8)) Or8_64 (.in0(wire_415), .in1({{7{1'b0}}, wire_341 }), .out(wire_201));
  TC_Constant # (.UUID(64'd378759622486388439 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFF006301)) Constant64_65 (.out(wire_338));
  TC_Constant # (.UUID(64'd4312411360349976773 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFF0002FF)) Constant64_66 (.out(wire_346));
  TC_LessU # (.UUID(64'd3095779165657668680 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_67 (.in0(wire_346), .in1(wire_62), .out(wire_287));
  TC_LessU # (.UUID(64'd1791836493397789689 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_68 (.in0(wire_62), .in1(wire_338), .out(wire_189));
  TC_And # (.UUID(64'd2636987386574953250 ^ UUID), .BIT_WIDTH(64'd1)) And_69 (.in0(wire_287), .in1(wire_189), .out(wire_403));
  TC_Shr # (.UUID(64'd3207325135725610088 ^ UUID), .BIT_WIDTH(64'd64)) Shr64_70 (.in(wire_62), .shift(wire_431), .out(wire_411));
  TC_Constant # (.UUID(64'd3459684029060330791 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_71 (.out(wire_431));
  TC_Add # (.UUID(64'd2236239263451235497 ^ UUID), .BIT_WIDTH(64'd64)) Add64_72 (.in0(wire_411), .in1(wire_383), .ci(1'd0), .out(wire_100), .co());
  TC_Constant # (.UUID(64'd1626638495718484720 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFC03FFF40)) Constant64_73 (.out(wire_383));
  TC_DotMatrixDisplay # (.UUID(64'd4245692389190270041 ^ UUID)) DotMatrixDisplay_74 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_26[0:0]), .color_info(wire_14), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1081087944869677309 ^ UUID)) DotMatrixDisplay_75 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_26[0:0]), .color_info(wire_106), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2014305234788474288 ^ UUID)) DotMatrixDisplay_76 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_26[0:0]), .color_info(wire_52), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1250514568413918296 ^ UUID)) DotMatrixDisplay_77 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_26[0:0]), .color_info(wire_58), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd4061792430659240502 ^ UUID)) DotMatrixDisplay_78 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_26[0:0]), .color_info(wire_23), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd3071246575142680608 ^ UUID)) DotMatrixDisplay_79 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_26[0:0]), .color_info(wire_68), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd3295334999887271511 ^ UUID)) DotMatrixDisplay_80 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_26[0:0]), .color_info(wire_79), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1871017718047496943 ^ UUID)) DotMatrixDisplay_81 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_26[0:0]), .color_info(wire_38), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2664915947813833550 ^ UUID)) DotMatrixDisplay_82 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_26[0:0]), .color_info(wire_55), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd3825264023869012084 ^ UUID)) DotMatrixDisplay_83 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_26[0:0]), .color_info(wire_10), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd629835669602455866 ^ UUID)) DotMatrixDisplay_84 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_26[0:0]), .color_info(wire_86), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd847161699868994951 ^ UUID)) DotMatrixDisplay_85 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_26[0:0]), .color_info(wire_76), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2130616956542995063 ^ UUID)) DotMatrixDisplay_86 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_26[0:0]), .color_info(wire_85), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd2711165688276813194 ^ UUID)) DotMatrixDisplay_87 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_26[0:0]), .color_info(wire_34), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1269560416894204461 ^ UUID)) DotMatrixDisplay_88 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_26[0:0]), .color_info(wire_22), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd3526909426203271252 ^ UUID)) DotMatrixDisplay_89 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_26[0:0]), .color_info(wire_39), .pixel_info(wire_26));
  TC_DotMatrixDisplay # (.UUID(64'd1847294820130042127 ^ UUID)) DotMatrixDisplay_90 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_24[0:0]), .color_info(wire_14), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd199253922724809882 ^ UUID)) DotMatrixDisplay_91 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_24[0:0]), .color_info(wire_106), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1667339508018048744 ^ UUID)) DotMatrixDisplay_92 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_24[0:0]), .color_info(wire_52), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1872596990519231642 ^ UUID)) DotMatrixDisplay_93 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_24[0:0]), .color_info(wire_58), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd3762393731378683491 ^ UUID)) DotMatrixDisplay_94 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_24[0:0]), .color_info(wire_23), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd3447451469009434368 ^ UUID)) DotMatrixDisplay_95 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_24[0:0]), .color_info(wire_68), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1557597890283114420 ^ UUID)) DotMatrixDisplay_96 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_24[0:0]), .color_info(wire_79), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1741251584214982772 ^ UUID)) DotMatrixDisplay_97 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_24[0:0]), .color_info(wire_38), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1378104951951587866 ^ UUID)) DotMatrixDisplay_98 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_24[0:0]), .color_info(wire_55), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd4173621311689271022 ^ UUID)) DotMatrixDisplay_99 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_24[0:0]), .color_info(wire_10), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd430601579600007200 ^ UUID)) DotMatrixDisplay_100 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_24[0:0]), .color_info(wire_86), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd2254006063250506991 ^ UUID)) DotMatrixDisplay_101 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_24[0:0]), .color_info(wire_76), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1888159867266837123 ^ UUID)) DotMatrixDisplay_102 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_24[0:0]), .color_info(wire_85), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1958363186366712055 ^ UUID)) DotMatrixDisplay_103 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_24[0:0]), .color_info(wire_34), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd2041128009341724824 ^ UUID)) DotMatrixDisplay_104 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_24[0:0]), .color_info(wire_22), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd3382347561032158534 ^ UUID)) DotMatrixDisplay_105 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_24[0:0]), .color_info(wire_39), .pixel_info(wire_24));
  TC_DotMatrixDisplay # (.UUID(64'd1602173510156883661 ^ UUID)) DotMatrixDisplay_106 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_42[0:0]), .color_info(wire_14), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1558734432975654504 ^ UUID)) DotMatrixDisplay_107 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_42[0:0]), .color_info(wire_106), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1844899675411949500 ^ UUID)) DotMatrixDisplay_108 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_42[0:0]), .color_info(wire_52), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd2753421226125773168 ^ UUID)) DotMatrixDisplay_109 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_42[0:0]), .color_info(wire_58), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1043017127660876480 ^ UUID)) DotMatrixDisplay_110 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_42[0:0]), .color_info(wire_23), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd2598571183317024345 ^ UUID)) DotMatrixDisplay_111 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_42[0:0]), .color_info(wire_68), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd807767532488760335 ^ UUID)) DotMatrixDisplay_112 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_42[0:0]), .color_info(wire_79), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1328285229437952766 ^ UUID)) DotMatrixDisplay_113 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_42[0:0]), .color_info(wire_38), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1078419801499832407 ^ UUID)) DotMatrixDisplay_114 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_42[0:0]), .color_info(wire_55), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1384507883605792292 ^ UUID)) DotMatrixDisplay_115 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_42[0:0]), .color_info(wire_10), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd491542944227860794 ^ UUID)) DotMatrixDisplay_116 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_42[0:0]), .color_info(wire_86), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd4013440861536287816 ^ UUID)) DotMatrixDisplay_117 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_42[0:0]), .color_info(wire_76), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1345021795193577811 ^ UUID)) DotMatrixDisplay_118 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_42[0:0]), .color_info(wire_85), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd3448147012112863839 ^ UUID)) DotMatrixDisplay_119 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_42[0:0]), .color_info(wire_34), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd3991347083632783865 ^ UUID)) DotMatrixDisplay_120 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_42[0:0]), .color_info(wire_22), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd1438929833035091957 ^ UUID)) DotMatrixDisplay_121 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_42[0:0]), .color_info(wire_39), .pixel_info(wire_42));
  TC_DotMatrixDisplay # (.UUID(64'd3507520420270208770 ^ UUID)) DotMatrixDisplay_122 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_44[0:0]), .color_info(wire_14), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1784882512189347093 ^ UUID)) DotMatrixDisplay_123 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_44[0:0]), .color_info(wire_106), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd2122312382829692208 ^ UUID)) DotMatrixDisplay_124 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_44[0:0]), .color_info(wire_52), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3141905182129353877 ^ UUID)) DotMatrixDisplay_125 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_44[0:0]), .color_info(wire_58), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3473597012091497710 ^ UUID)) DotMatrixDisplay_126 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_44[0:0]), .color_info(wire_23), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1808490368191185449 ^ UUID)) DotMatrixDisplay_127 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_44[0:0]), .color_info(wire_68), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1562987427505910492 ^ UUID)) DotMatrixDisplay_128 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_44[0:0]), .color_info(wire_79), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1963694696365273293 ^ UUID)) DotMatrixDisplay_129 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_44[0:0]), .color_info(wire_38), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3452649505164889566 ^ UUID)) DotMatrixDisplay_130 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_44[0:0]), .color_info(wire_55), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd4074866046846024365 ^ UUID)) DotMatrixDisplay_131 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_44[0:0]), .color_info(wire_10), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3421062344287591638 ^ UUID)) DotMatrixDisplay_132 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_44[0:0]), .color_info(wire_86), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1656817259187101187 ^ UUID)) DotMatrixDisplay_133 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_44[0:0]), .color_info(wire_76), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1828136908011057645 ^ UUID)) DotMatrixDisplay_134 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_44[0:0]), .color_info(wire_85), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3938622764814591470 ^ UUID)) DotMatrixDisplay_135 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_44[0:0]), .color_info(wire_34), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3977226084215625849 ^ UUID)) DotMatrixDisplay_136 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_44[0:0]), .color_info(wire_22), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd3624336617201189335 ^ UUID)) DotMatrixDisplay_137 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_44[0:0]), .color_info(wire_39), .pixel_info(wire_44));
  TC_DotMatrixDisplay # (.UUID(64'd1051202942619435355 ^ UUID)) DotMatrixDisplay_138 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_2[0:0]), .color_info(wire_14), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1155289762323060933 ^ UUID)) DotMatrixDisplay_139 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_2[0:0]), .color_info(wire_106), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd4519341567349756337 ^ UUID)) DotMatrixDisplay_140 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_2[0:0]), .color_info(wire_52), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2722966304414546736 ^ UUID)) DotMatrixDisplay_141 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_2[0:0]), .color_info(wire_58), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd209028992023888191 ^ UUID)) DotMatrixDisplay_142 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_2[0:0]), .color_info(wire_23), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1240341250017908700 ^ UUID)) DotMatrixDisplay_143 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_2[0:0]), .color_info(wire_68), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3929540560851822745 ^ UUID)) DotMatrixDisplay_144 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_2[0:0]), .color_info(wire_79), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3966679511028762021 ^ UUID)) DotMatrixDisplay_145 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_2[0:0]), .color_info(wire_38), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd69502193858986266 ^ UUID)) DotMatrixDisplay_146 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_2[0:0]), .color_info(wire_55), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd41038936696827963 ^ UUID)) DotMatrixDisplay_147 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_2[0:0]), .color_info(wire_10), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2054359701663655273 ^ UUID)) DotMatrixDisplay_148 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_2[0:0]), .color_info(wire_86), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd2424292374505990024 ^ UUID)) DotMatrixDisplay_149 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_2[0:0]), .color_info(wire_76), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1922480469082329831 ^ UUID)) DotMatrixDisplay_150 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_2[0:0]), .color_info(wire_85), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3477201688326722707 ^ UUID)) DotMatrixDisplay_151 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_2[0:0]), .color_info(wire_34), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd3497841040434478899 ^ UUID)) DotMatrixDisplay_152 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_2[0:0]), .color_info(wire_22), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1983868183368881738 ^ UUID)) DotMatrixDisplay_153 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_2[0:0]), .color_info(wire_39), .pixel_info(wire_2));
  TC_DotMatrixDisplay # (.UUID(64'd1429891968970895491 ^ UUID)) DotMatrixDisplay_154 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_30[0:0]), .color_info(wire_14), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd143829235001463726 ^ UUID)) DotMatrixDisplay_155 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_30[0:0]), .color_info(wire_106), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd112444896658137125 ^ UUID)) DotMatrixDisplay_156 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_30[0:0]), .color_info(wire_52), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2701201058716092627 ^ UUID)) DotMatrixDisplay_157 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_30[0:0]), .color_info(wire_58), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd1729038379468812768 ^ UUID)) DotMatrixDisplay_158 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_30[0:0]), .color_info(wire_23), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd94168968341889190 ^ UUID)) DotMatrixDisplay_159 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_30[0:0]), .color_info(wire_68), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2683831824093842119 ^ UUID)) DotMatrixDisplay_160 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_30[0:0]), .color_info(wire_79), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2426582617545712316 ^ UUID)) DotMatrixDisplay_161 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_30[0:0]), .color_info(wire_38), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd703010574784385063 ^ UUID)) DotMatrixDisplay_162 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_30[0:0]), .color_info(wire_55), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd4494316196581305812 ^ UUID)) DotMatrixDisplay_163 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_30[0:0]), .color_info(wire_10), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3916490575512509304 ^ UUID)) DotMatrixDisplay_164 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_30[0:0]), .color_info(wire_86), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2751814764301207852 ^ UUID)) DotMatrixDisplay_165 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_30[0:0]), .color_info(wire_76), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd4469838669328512932 ^ UUID)) DotMatrixDisplay_166 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_30[0:0]), .color_info(wire_85), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3408293338592194612 ^ UUID)) DotMatrixDisplay_167 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_30[0:0]), .color_info(wire_34), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd199805756176147134 ^ UUID)) DotMatrixDisplay_168 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_30[0:0]), .color_info(wire_22), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd2141840590039932523 ^ UUID)) DotMatrixDisplay_169 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_30[0:0]), .color_info(wire_39), .pixel_info(wire_30));
  TC_DotMatrixDisplay # (.UUID(64'd3855379692753837257 ^ UUID)) DotMatrixDisplay_170 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_104[0:0]), .color_info(wire_14), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd2531282466371223794 ^ UUID)) DotMatrixDisplay_171 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_104[0:0]), .color_info(wire_106), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd3266338675676829761 ^ UUID)) DotMatrixDisplay_172 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_104[0:0]), .color_info(wire_52), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd4389367126554349096 ^ UUID)) DotMatrixDisplay_173 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_104[0:0]), .color_info(wire_58), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd4464643644768383458 ^ UUID)) DotMatrixDisplay_174 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_104[0:0]), .color_info(wire_23), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd2316679577792341300 ^ UUID)) DotMatrixDisplay_175 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_104[0:0]), .color_info(wire_68), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd1284989749365717974 ^ UUID)) DotMatrixDisplay_176 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_104[0:0]), .color_info(wire_79), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd3358879124586778308 ^ UUID)) DotMatrixDisplay_177 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_104[0:0]), .color_info(wire_38), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd3892470599579388761 ^ UUID)) DotMatrixDisplay_178 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_104[0:0]), .color_info(wire_55), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd2409555869879819577 ^ UUID)) DotMatrixDisplay_179 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_104[0:0]), .color_info(wire_10), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd2470242801042046595 ^ UUID)) DotMatrixDisplay_180 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_104[0:0]), .color_info(wire_86), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd4444749580746722924 ^ UUID)) DotMatrixDisplay_181 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_104[0:0]), .color_info(wire_76), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd2244020422625260257 ^ UUID)) DotMatrixDisplay_182 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_104[0:0]), .color_info(wire_85), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd3298188220166804620 ^ UUID)) DotMatrixDisplay_183 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_104[0:0]), .color_info(wire_34), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd137780235944102946 ^ UUID)) DotMatrixDisplay_184 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_104[0:0]), .color_info(wire_22), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd346284501654386559 ^ UUID)) DotMatrixDisplay_185 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_104[0:0]), .color_info(wire_39), .pixel_info(wire_104));
  TC_DotMatrixDisplay # (.UUID(64'd114465287468131338 ^ UUID)) DotMatrixDisplay_186 (.clk(clk), .rst(rst), .en_y(wire_14[0:0]), .en_x(wire_91[0:0]), .color_info(wire_14), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd527271392111862154 ^ UUID)) DotMatrixDisplay_187 (.clk(clk), .rst(rst), .en_y(wire_106[0:0]), .en_x(wire_91[0:0]), .color_info(wire_106), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd1364848831498191197 ^ UUID)) DotMatrixDisplay_188 (.clk(clk), .rst(rst), .en_y(wire_52[0:0]), .en_x(wire_91[0:0]), .color_info(wire_52), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd1949485794081205826 ^ UUID)) DotMatrixDisplay_189 (.clk(clk), .rst(rst), .en_y(wire_58[0:0]), .en_x(wire_91[0:0]), .color_info(wire_58), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd1516290122148093922 ^ UUID)) DotMatrixDisplay_190 (.clk(clk), .rst(rst), .en_y(wire_23[0:0]), .en_x(wire_91[0:0]), .color_info(wire_23), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd1208061358446223542 ^ UUID)) DotMatrixDisplay_191 (.clk(clk), .rst(rst), .en_y(wire_68[0:0]), .en_x(wire_91[0:0]), .color_info(wire_68), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd1801161967132270202 ^ UUID)) DotMatrixDisplay_192 (.clk(clk), .rst(rst), .en_y(wire_79[0:0]), .en_x(wire_91[0:0]), .color_info(wire_79), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd2045142587737685395 ^ UUID)) DotMatrixDisplay_193 (.clk(clk), .rst(rst), .en_y(wire_38[0:0]), .en_x(wire_91[0:0]), .color_info(wire_38), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd2448973839005186099 ^ UUID)) DotMatrixDisplay_194 (.clk(clk), .rst(rst), .en_y(wire_55[0:0]), .en_x(wire_91[0:0]), .color_info(wire_55), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd3541848710978226558 ^ UUID)) DotMatrixDisplay_195 (.clk(clk), .rst(rst), .en_y(wire_10[0:0]), .en_x(wire_91[0:0]), .color_info(wire_10), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd4052483778756570721 ^ UUID)) DotMatrixDisplay_196 (.clk(clk), .rst(rst), .en_y(wire_86[0:0]), .en_x(wire_91[0:0]), .color_info(wire_86), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd3617339000090961038 ^ UUID)) DotMatrixDisplay_197 (.clk(clk), .rst(rst), .en_y(wire_76[0:0]), .en_x(wire_91[0:0]), .color_info(wire_76), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd870007035309902639 ^ UUID)) DotMatrixDisplay_198 (.clk(clk), .rst(rst), .en_y(wire_85[0:0]), .en_x(wire_91[0:0]), .color_info(wire_85), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd2064733774029395729 ^ UUID)) DotMatrixDisplay_199 (.clk(clk), .rst(rst), .en_y(wire_34[0:0]), .en_x(wire_91[0:0]), .color_info(wire_34), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd2409151620052632979 ^ UUID)) DotMatrixDisplay_200 (.clk(clk), .rst(rst), .en_y(wire_22[0:0]), .en_x(wire_91[0:0]), .color_info(wire_22), .pixel_info(wire_91));
  TC_DotMatrixDisplay # (.UUID(64'd3264256391491672189 ^ UUID)) DotMatrixDisplay_201 (.clk(clk), .rst(rst), .en_y(wire_39[0:0]), .en_x(wire_91[0:0]), .color_info(wire_39), .pixel_info(wire_91));
  Instructionz_Decoder # (.UUID(64'd2879907105418065125 ^ UUID)) Instructionz_Decoder_202 (.clk(clk), .rst(rst), .Input(wire_243), .Enabled(wire_261), .ALU(wire_90), .Control(wire_93), .Memory_Read(wire_141), .Fence(wire_418), .System(wire_237), .Error(wire_384));
  Programz_Counter # (.UUID(64'd4003924343034246755 ^ UUID)) Programz_Counter_203 (.clk(clk), .rst(rst), .Input(wire_325), .Override(wire_281), .Enable(wire_373), .Value(wire_227), .Output(wire_105));
  Controlz_Block # (.UUID(64'd3143867639452171112 ^ UUID)) Controlz_Block_204 (.clk(clk), .rst(rst), .Instruction(wire_243), .Register_1(wire_15), .Register_2(wire_256), .Enabled(wire_93), .PC(wire_105), .Register_Out(wire_1_1), .Write_Register(wire_157), .PC_Out(wire_227), .Should_Jump(wire_281));
  ALU # (.UUID(64'd2776056562894842104 ^ UUID)) ALU_205 (.clk(clk), .rst(rst), .Register_1(wire_15), .Register_2(wire_256), .Instruction(wire_243), .Enable(wire_90), .PC(wire_105), .Error(wire_395), .Output(wire_1_0));
  Displayz_Controller # (.UUID(64'd2341064131763610923 ^ UUID)) Displayz_Controller_206 (.clk(clk), .rst(rst), .Value(wire_9[31:0]), .Enable(wire_403), .Address(wire_100[31:0]), .Output_1(wire_14), .Output_2(wire_106), .Output_3(wire_52), .Output_4(wire_58), .Output_5(wire_23), .Output_6(wire_68), .Output_7(wire_79), .Output_8(wire_38), .Output_9(wire_55), .Output_10(wire_10), .Output_11(wire_86), .Output_12(wire_76), .Output_13(wire_85), .Output_14(wire_34), .Output_15(wire_22), .Output_16(wire_39), .Output_17(wire_26), .Output_18(wire_24), .Output_19(wire_42), .Output_20(wire_44), .Output_21(wire_2), .Output_22(wire_30), .Output_23(wire_104), .Output_24(wire_91));
  TC_Splitter32 # (.UUID(64'd2772194238259801067 ^ UUID)) Splitter32_207 (.in(wire_322), .out0(wire_321), .out1(wire_82), .out2(), .out3());
  TC_Switch # (.UUID(64'd3249943738321454775 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_208 (.en(wire_355), .in(wire_137), .out(wire_322));
  TC_Splitter8 # (.UUID(64'd1406322775684055465 ^ UUID)) Splitter8_209 (.in(wire_321), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_288));
  TC_Splitter8 # (.UUID(64'd2176169810335608793 ^ UUID)) Splitter8_210 (.in(wire_82), .out0(wire_340), .out1(wire_102), .out2(wire_195), .out3(wire_71), .out4(), .out5(), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd2122703970950031676 ^ UUID)) Splitter32_211 (.in(wire_137), .out0(), .out1(wire_275), .out2(wire_318), .out3());
  TC_Splitter8 # (.UUID(64'd2766344383163818103 ^ UUID)) Splitter8_212 (.in(wire_275), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_84));
  TC_Splitter8 # (.UUID(64'd693403901791489341 ^ UUID)) Splitter8_213 (.in(wire_318), .out0(wire_332), .out1(wire_220), .out2(wire_301), .out3(wire_449), .out4(), .out5(), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd2382784469017292456 ^ UUID)) Splitter32_214 (.in(wire_137), .out0(), .out1(), .out2(wire_316), .out3(wire_298));
  TC_Splitter8 # (.UUID(64'd1544065967333299809 ^ UUID)) Splitter8_215 (.in(wire_316), .out0(), .out1(), .out2(), .out3(), .out4(wire_364), .out5(wire_382), .out6(wire_158), .out7(wire_343));
  TC_Splitter8 # (.UUID(64'd3539257858633878690 ^ UUID)) Splitter8_216 (.in(wire_298), .out0(wire_363), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Register # (.UUID(64'd2434775662967180197 ^ UUID), .BIT_WIDTH(64'd32)) Register32_217 (.clk(clk), .rst(rst), .load(wire_442), .save(wire_312), .in(wire_1), .out(wire_53));
  TC_Constant # (.UUID(64'd1802124805265315764 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_218 (.out(wire_442));
  TC_Register # (.UUID(64'd1476595443994256450 ^ UUID), .BIT_WIDTH(64'd32)) Register32_219 (.clk(clk), .rst(rst), .load(wire_302), .save(wire_194), .in(wire_1), .out(wire_214));
  TC_Constant # (.UUID(64'd906466517651869234 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_220 (.out(wire_302));
  TC_Register # (.UUID(64'd2873357547679377394 ^ UUID), .BIT_WIDTH(64'd32)) Register32_221 (.clk(clk), .rst(rst), .load(wire_412), .save(wire_239), .in(wire_1), .out(wire_176));
  TC_Constant # (.UUID(64'd3666464021175878387 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_222 (.out(wire_412));
  TC_Register # (.UUID(64'd561277027413541936 ^ UUID), .BIT_WIDTH(64'd32)) Register32_223 (.clk(clk), .rst(rst), .load(wire_420), .save(wire_225), .in(wire_1), .out(wire_135));
  TC_Constant # (.UUID(64'd4050205726037109794 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_224 (.out(wire_420));
  TC_Register # (.UUID(64'd3403507603070574860 ^ UUID), .BIT_WIDTH(64'd32)) Register32_225 (.clk(clk), .rst(rst), .load(wire_83), .save(wire_352), .in(wire_1), .out(wire_118));
  TC_Constant # (.UUID(64'd2178507116231302121 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_226 (.out(wire_83));
  TC_Register # (.UUID(64'd1426880244683972691 ^ UUID), .BIT_WIDTH(64'd32)) Register32_227 (.clk(clk), .rst(rst), .load(wire_207), .save(wire_271), .in(wire_1), .out(wire_173));
  TC_Constant # (.UUID(64'd3825326989900596455 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_228 (.out(wire_207));
  TC_Register # (.UUID(64'd1433639157801468264 ^ UUID), .BIT_WIDTH(64'd32)) Register32_229 (.clk(clk), .rst(rst), .load(wire_178), .save(wire_428), .in(wire_1), .out(wire_45));
  TC_Constant # (.UUID(64'd292725899645715216 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_230 (.out(wire_178));
  TC_Splitter8 # (.UUID(64'd1653133521485656185 ^ UUID)) Splitter8_231 (.in(wire_274), .out0(), .out1(wire_312), .out2(wire_194), .out3(wire_239), .out4(wire_225), .out5(wire_352), .out6(wire_271), .out7(wire_428));
  TC_Splitter32 # (.UUID(64'd1690400056863910564 ^ UUID)) Splitter32_232 (.in(wire_78), .out0(wire_274), .out1(wire_148), .out2(wire_32), .out3(wire_216));
  TC_Register # (.UUID(64'd2143354438073683198 ^ UUID), .BIT_WIDTH(64'd32)) Register32_233 (.clk(clk), .rst(rst), .load(wire_327), .save(wire_375), .in(wire_1), .out(wire_215));
  TC_Constant # (.UUID(64'd436819717719264517 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_234 (.out(wire_327));
  TC_Register # (.UUID(64'd2590062290789180301 ^ UUID), .BIT_WIDTH(64'd32)) Register32_235 (.clk(clk), .rst(rst), .load(wire_196), .save(wire_278), .in(wire_1), .out(wire_162));
  TC_Constant # (.UUID(64'd2714367564197902483 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_236 (.out(wire_196));
  TC_Register # (.UUID(64'd1660484509566904138 ^ UUID), .BIT_WIDTH(64'd32)) Register32_237 (.clk(clk), .rst(rst), .load(wire_334), .save(wire_270), .in(wire_1), .out(wire_116));
  TC_Constant # (.UUID(64'd1855739425211009605 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_238 (.out(wire_334));
  TC_Register # (.UUID(64'd2903681585765584581 ^ UUID), .BIT_WIDTH(64'd32)) Register32_239 (.clk(clk), .rst(rst), .load(wire_447), .save(wire_50), .in(wire_1), .out(wire_126));
  TC_Constant # (.UUID(64'd3943230229408446956 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_240 (.out(wire_447));
  TC_Register # (.UUID(64'd1154702339103748081 ^ UUID), .BIT_WIDTH(64'd32)) Register32_241 (.clk(clk), .rst(rst), .load(wire_308), .save(wire_120), .in(wire_1), .out(wire_198));
  TC_Constant # (.UUID(64'd2782535415991006015 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_242 (.out(wire_308));
  TC_Register # (.UUID(64'd3879850639627936494 ^ UUID), .BIT_WIDTH(64'd32)) Register32_243 (.clk(clk), .rst(rst), .load(wire_401), .save(wire_361), .in(wire_1), .out(wire_88));
  TC_Constant # (.UUID(64'd3274576321670644412 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_244 (.out(wire_401));
  TC_Register # (.UUID(64'd750146477149948725 ^ UUID), .BIT_WIDTH(64'd32)) Register32_245 (.clk(clk), .rst(rst), .load(wire_446), .save(wire_354), .in(wire_1), .out(wire_228));
  TC_Constant # (.UUID(64'd4179987660858840768 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_246 (.out(wire_446));
  TC_Register # (.UUID(64'd3839315151889669018 ^ UUID), .BIT_WIDTH(64'd32)) Register32_247 (.clk(clk), .rst(rst), .load(wire_357), .save(wire_49), .in(wire_1), .out(wire_111));
  TC_Constant # (.UUID(64'd3591114557495138038 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_248 (.out(wire_357));
  TC_Splitter8 # (.UUID(64'd4499458438455487445 ^ UUID)) Splitter8_249 (.in(wire_148), .out0(wire_375), .out1(wire_278), .out2(wire_270), .out3(wire_50), .out4(wire_120), .out5(wire_361), .out6(wire_354), .out7(wire_49));
  TC_Register # (.UUID(64'd2699651052599423094 ^ UUID), .BIT_WIDTH(64'd32)) Register32_250 (.clk(clk), .rst(rst), .load(wire_405), .save(wire_138), .in(wire_1), .out(wire_99));
  TC_Constant # (.UUID(64'd825394209917224559 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_251 (.out(wire_405));
  TC_Register # (.UUID(64'd4384947640070513041 ^ UUID), .BIT_WIDTH(64'd32)) Register32_252 (.clk(clk), .rst(rst), .load(wire_61), .save(wire_16), .in(wire_1), .out(wire_63));
  TC_Constant # (.UUID(64'd784266035874962889 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_253 (.out(wire_61));
  TC_Register # (.UUID(64'd2229426681918121128 ^ UUID), .BIT_WIDTH(64'd32)) Register32_254 (.clk(clk), .rst(rst), .load(wire_410), .save(wire_101), .in(wire_1), .out(wire_267));
  TC_Constant # (.UUID(64'd152278999248324997 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_255 (.out(wire_410));
  TC_Register # (.UUID(64'd3268871637652075343 ^ UUID), .BIT_WIDTH(64'd32)) Register32_256 (.clk(clk), .rst(rst), .load(wire_177), .save(wire_161), .in(wire_1), .out(wire_95));
  TC_Constant # (.UUID(64'd1908821689548691242 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_257 (.out(wire_177));
  TC_Register # (.UUID(64'd1970684396627040945 ^ UUID), .BIT_WIDTH(64'd32)) Register32_258 (.clk(clk), .rst(rst), .load(wire_236), .save(wire_139), .in(wire_1), .out(wire_179));
  TC_Constant # (.UUID(64'd4480038280979685486 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_259 (.out(wire_236));
  TC_Register # (.UUID(64'd3497136520650075956 ^ UUID), .BIT_WIDTH(64'd32)) Register32_260 (.clk(clk), .rst(rst), .load(wire_259), .save(wire_235), .in(wire_1), .out(wire_21));
  TC_Constant # (.UUID(64'd1621579246550563398 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_261 (.out(wire_259));
  TC_Register # (.UUID(64'd1237076464754429007 ^ UUID), .BIT_WIDTH(64'd32)) Register32_262 (.clk(clk), .rst(rst), .load(wire_390), .save(wire_132), .in(wire_1), .out(wire_128));
  TC_Constant # (.UUID(64'd2701540367966331248 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_263 (.out(wire_390));
  TC_Register # (.UUID(64'd1951931176718714339 ^ UUID), .BIT_WIDTH(64'd32)) Register32_264 (.clk(clk), .rst(rst), .load(wire_417), .save(wire_47), .in(wire_1), .out(wire_159));
  TC_Constant # (.UUID(64'd3413647735577703717 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_265 (.out(wire_417));
  TC_Splitter8 # (.UUID(64'd1256689854284230608 ^ UUID)) Splitter8_266 (.in(wire_32), .out0(wire_138), .out1(wire_16), .out2(wire_101), .out3(wire_161), .out4(wire_139), .out5(wire_235), .out6(wire_132), .out7(wire_47));
  TC_Register # (.UUID(64'd1202578987467448203 ^ UUID), .BIT_WIDTH(64'd32)) Register32_267 (.clk(clk), .rst(rst), .load(wire_377), .save(wire_263), .in(wire_1), .out(wire_110));
  TC_Constant # (.UUID(64'd1548053689714413518 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_268 (.out(wire_377));
  TC_Register # (.UUID(64'd4537541985681412933 ^ UUID), .BIT_WIDTH(64'd32)) Register32_269 (.clk(clk), .rst(rst), .load(wire_407), .save(wire_234), .in(wire_1), .out(wire_249));
  TC_Constant # (.UUID(64'd2882491480880030580 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_270 (.out(wire_407));
  TC_Register # (.UUID(64'd3004932813165070893 ^ UUID), .BIT_WIDTH(64'd32)) Register32_271 (.clk(clk), .rst(rst), .load(wire_397), .save(wire_57), .in(wire_1), .out(wire_28));
  TC_Constant # (.UUID(64'd1225443957963169271 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_272 (.out(wire_397));
  TC_Register # (.UUID(64'd1678989197830856400 ^ UUID), .BIT_WIDTH(64'd32)) Register32_273 (.clk(clk), .rst(rst), .load(wire_404), .save(wire_244), .in(wire_1), .out(wire_37));
  TC_Constant # (.UUID(64'd1594982685616301849 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_274 (.out(wire_404));
  TC_Register # (.UUID(64'd1577322723702123335 ^ UUID), .BIT_WIDTH(64'd32)) Register32_275 (.clk(clk), .rst(rst), .load(wire_387), .save(wire_35), .in(wire_1), .out(wire_96));
  TC_Constant # (.UUID(64'd3887081089242553540 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_276 (.out(wire_387));
  TC_Register # (.UUID(64'd755291711939798802 ^ UUID), .BIT_WIDTH(64'd32)) Register32_277 (.clk(clk), .rst(rst), .load(wire_92), .save(wire_202), .in(wire_1), .out(wire_3));
  TC_Constant # (.UUID(64'd2103787712320682162 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_278 (.out(wire_92));
  TC_Register # (.UUID(64'd1800689002083486681 ^ UUID), .BIT_WIDTH(64'd32)) Register32_279 (.clk(clk), .rst(rst), .load(wire_413), .save(wire_229), .in(wire_1), .out(wire_150));
  TC_Constant # (.UUID(64'd2511022624567749327 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_280 (.out(wire_413));
  TC_Register # (.UUID(64'd994756424935798740 ^ UUID), .BIT_WIDTH(64'd32)) Register32_281 (.clk(clk), .rst(rst), .load(wire_358), .save(wire_282), .in(wire_1), .out(wire_221));
  TC_Constant # (.UUID(64'd2795214332012202500 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_282 (.out(wire_358));
  TC_Splitter8 # (.UUID(64'd1416078167936227239 ^ UUID)) Splitter8_283 (.in(wire_216), .out0(wire_263), .out1(wire_234), .out2(wire_57), .out3(wire_244), .out4(wire_35), .out5(wire_202), .out6(wire_229), .out7(wire_282));
  TC_Buffer # (.UUID(64'd2795247990498223635 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_284 (.in(wire_243), .out(wire_137));
  TC_Switch # (.UUID(64'd2309169332765144302 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_285 (.en(wire_77), .in(wire_311), .out(wire_167_4));
  TC_Switch # (.UUID(64'd4273634959314961929 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_286 (.en(wire_27), .in(wire_53), .out(wire_167_2));
  TC_Switch # (.UUID(64'd4067802285386255953 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_287 (.en(wire_266), .in(wire_214), .out(wire_167_0));
  TC_Switch # (.UUID(64'd1273525424053278178 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_288 (.en(wire_262), .in(wire_176), .out(wire_167_1));
  TC_Switch # (.UUID(64'd3315808851101833106 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_289 (.en(wire_253), .in(wire_135), .out(wire_167_3));
  TC_Switch # (.UUID(64'd4398866812963762499 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_290 (.en(wire_170), .in(wire_118), .out(wire_167_5));
  TC_Switch # (.UUID(64'd1809351694222139092 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_291 (.en(wire_124), .in(wire_173), .out(wire_167_6));
  TC_Switch # (.UUID(64'd1083920152741857132 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_292 (.en(wire_59), .in(wire_45), .out(wire_167_7));
  TC_Splitter8 # (.UUID(64'd651420256423447480 ^ UUID)) Splitter8_293 (.in(wire_331), .out0(wire_77), .out1(wire_27), .out2(wire_266), .out3(wire_262), .out4(wire_253), .out5(wire_170), .out6(wire_124), .out7(wire_59));
  TC_Splitter32 # (.UUID(64'd2226110187981876694 ^ UUID)) Splitter32_294 (.in(wire_315), .out0(wire_331), .out1(wire_72), .out2(wire_277), .out3(wire_213));
  TC_Switch # (.UUID(64'd2766902449608102218 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_295 (.en(wire_223), .in(wire_311), .out(wire_70_8));
  TC_Switch # (.UUID(64'd2860593462451573679 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_296 (.en(wire_54), .in(wire_53), .out(wire_70_6));
  TC_Switch # (.UUID(64'd4428495750854660128 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_297 (.en(wire_200), .in(wire_214), .out(wire_70_4));
  TC_Switch # (.UUID(64'd4465516763146188498 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_298 (.en(wire_204), .in(wire_176), .out(wire_70_2));
  TC_Switch # (.UUID(64'd3599770261062141485 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_299 (.en(wire_152), .in(wire_135), .out(wire_70_0));
  TC_Switch # (.UUID(64'd1576641770439589705 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_300 (.en(wire_127), .in(wire_118), .out(wire_70_1));
  TC_Switch # (.UUID(64'd3557889408083951009 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_301 (.en(wire_238), .in(wire_173), .out(wire_70_3));
  TC_Switch # (.UUID(64'd297128742924195800 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_302 (.en(wire_140), .in(wire_45), .out(wire_70_5));
  TC_Splitter8 # (.UUID(64'd3661031462686444805 ^ UUID)) Splitter8_303 (.in(wire_51), .out0(wire_223), .out1(wire_54), .out2(wire_200), .out3(wire_204), .out4(wire_152), .out5(wire_127), .out6(wire_238), .out7(wire_140));
  TC_Splitter32 # (.UUID(64'd4478028120254975927 ^ UUID)) Splitter32_304 (.in(wire_432), .out0(wire_51), .out1(wire_319), .out2(wire_74), .out3(wire_199));
  TC_Switch # (.UUID(64'd2687210642419233272 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_305 (.en(wire_368), .in(wire_215), .out(wire_167_8));
  TC_Switch # (.UUID(64'd2642052529551879137 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_306 (.en(wire_381), .in(wire_162), .out(wire_167_9));
  TC_Switch # (.UUID(64'd2785323812348768480 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_307 (.en(wire_149), .in(wire_116), .out(wire_167_10));
  TC_Switch # (.UUID(64'd1116222274404407078 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_308 (.en(wire_230), .in(wire_126), .out(wire_167_11));
  TC_Switch # (.UUID(64'd398386866777763789 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_309 (.en(wire_103), .in(wire_198), .out(wire_167_12));
  TC_Switch # (.UUID(64'd1733035639828593569 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_310 (.en(wire_402), .in(wire_88), .out(wire_167_13));
  TC_Switch # (.UUID(64'd2051073364864718303 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_311 (.en(wire_134), .in(wire_228), .out(wire_167_14));
  TC_Switch # (.UUID(64'd330581453436973031 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_312 (.en(wire_423), .in(wire_111), .out(wire_167_15));
  TC_Splitter8 # (.UUID(64'd889672390800381668 ^ UUID)) Splitter8_313 (.in(wire_72), .out0(wire_368), .out1(wire_381), .out2(wire_149), .out3(wire_230), .out4(wire_103), .out5(wire_402), .out6(wire_134), .out7(wire_423));
  TC_Switch # (.UUID(64'd2661872456585422251 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_314 (.en(wire_206), .in(wire_215), .out(wire_70_7));
  TC_Switch # (.UUID(64'd1242802444509495187 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_315 (.en(wire_89), .in(wire_162), .out(wire_70_9));
  TC_Switch # (.UUID(64'd4222358155486673059 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_316 (.en(wire_240), .in(wire_116), .out(wire_70_10));
  TC_Switch # (.UUID(64'd2245412691587635604 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_317 (.en(wire_41), .in(wire_126), .out(wire_70_11));
  TC_Switch # (.UUID(64'd4125097606679472433 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_318 (.en(wire_303), .in(wire_198), .out(wire_70_12));
  TC_Switch # (.UUID(64'd1040059646614541790 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_319 (.en(wire_97), .in(wire_88), .out(wire_70_13));
  TC_Switch # (.UUID(64'd2616170767148541986 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_320 (.en(wire_276), .in(wire_228), .out(wire_70_14));
  TC_Switch # (.UUID(64'd862708665044883489 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_321 (.en(wire_374), .in(wire_111), .out(wire_70_15));
  TC_Splitter8 # (.UUID(64'd4406757921817552196 ^ UUID)) Splitter8_322 (.in(wire_319), .out0(wire_206), .out1(wire_89), .out2(wire_240), .out3(wire_41), .out4(wire_303), .out5(wire_97), .out6(wire_276), .out7(wire_374));
  TC_Switch # (.UUID(64'd2933115361403480394 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_323 (.en(wire_309), .in(wire_99), .out(wire_167_16));
  TC_Switch # (.UUID(64'd3666325126359315190 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_324 (.en(wire_219), .in(wire_63), .out(wire_167_17));
  TC_Switch # (.UUID(64'd3454177350459774129 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_325 (.en(wire_299), .in(wire_267), .out(wire_167_18));
  TC_Switch # (.UUID(64'd1302064961008901288 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_326 (.en(wire_398), .in(wire_95), .out(wire_167_19));
  TC_Switch # (.UUID(64'd3050102379920198435 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_327 (.en(wire_12), .in(wire_179), .out(wire_167_20));
  TC_Switch # (.UUID(64'd3248547773758430850 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_328 (.en(wire_426), .in(wire_21), .out(wire_167_21));
  TC_Switch # (.UUID(64'd2392548846227095871 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_329 (.en(wire_5), .in(wire_128), .out(wire_167_22));
  TC_Switch # (.UUID(64'd2108895439525214917 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_330 (.en(wire_290), .in(wire_159), .out(wire_167_23));
  TC_Splitter8 # (.UUID(64'd734113506290029937 ^ UUID)) Splitter8_331 (.in(wire_277), .out0(wire_309), .out1(wire_219), .out2(wire_299), .out3(wire_398), .out4(wire_12), .out5(wire_426), .out6(wire_5), .out7(wire_290));
  TC_Switch # (.UUID(64'd3661124640572735734 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_332 (.en(wire_183), .in(wire_99), .out(wire_70_16));
  TC_Switch # (.UUID(64'd3759680237115020462 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_333 (.en(wire_205), .in(wire_63), .out(wire_70_17));
  TC_Switch # (.UUID(64'd4381238231899394671 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_334 (.en(wire_289), .in(wire_267), .out(wire_70_18));
  TC_Switch # (.UUID(64'd4482953208222832838 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_335 (.en(wire_166), .in(wire_95), .out(wire_70_19));
  TC_Switch # (.UUID(64'd3776606891245099349 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_336 (.en(wire_347), .in(wire_179), .out(wire_70_20));
  TC_Switch # (.UUID(64'd2234887317273419702 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_337 (.en(wire_163), .in(wire_21), .out(wire_70_21));
  TC_Switch # (.UUID(64'd3003219917340010386 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_338 (.en(wire_80), .in(wire_128), .out(wire_70_22));
  TC_Switch # (.UUID(64'd3097210689935334749 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_339 (.en(wire_294), .in(wire_159), .out(wire_70_23));
  TC_Splitter8 # (.UUID(64'd366991715527825476 ^ UUID)) Splitter8_340 (.in(wire_74), .out0(wire_183), .out1(wire_205), .out2(wire_289), .out3(wire_166), .out4(wire_347), .out5(wire_163), .out6(wire_80), .out7(wire_294));
  TC_Switch # (.UUID(64'd3333625114167872620 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_341 (.en(wire_406), .in(wire_110), .out(wire_167_24));
  TC_Switch # (.UUID(64'd2355297711672223846 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_342 (.en(wire_248), .in(wire_249), .out(wire_167_25));
  TC_Switch # (.UUID(64'd592838331050856624 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_343 (.en(wire_112), .in(wire_28), .out(wire_167_26));
  TC_Switch # (.UUID(64'd3767868560430098562 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_344 (.en(wire_252), .in(wire_37), .out(wire_167_27));
  TC_Switch # (.UUID(64'd2192774683783783560 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_345 (.en(wire_292), .in(wire_96), .out(wire_167_28));
  TC_Switch # (.UUID(64'd670078746238553433 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_346 (.en(wire_94), .in(wire_3), .out(wire_167_29));
  TC_Switch # (.UUID(64'd3925537490124508737 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_347 (.en(wire_175), .in(wire_150), .out(wire_167_30));
  TC_Switch # (.UUID(64'd3338338420054904462 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_348 (.en(wire_250), .in(wire_221), .out(wire_167_31));
  TC_Splitter8 # (.UUID(64'd516961720266919740 ^ UUID)) Splitter8_349 (.in(wire_213), .out0(wire_406), .out1(wire_248), .out2(wire_112), .out3(wire_252), .out4(wire_292), .out5(wire_94), .out6(wire_175), .out7(wire_250));
  TC_Switch # (.UUID(64'd4574985456382582030 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_350 (.en(wire_188), .in(wire_110), .out(wire_70_24));
  TC_Switch # (.UUID(64'd2659320976288313996 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_351 (.en(wire_11), .in(wire_249), .out(wire_70_25));
  TC_Switch # (.UUID(64'd3224735037528383850 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_352 (.en(wire_122), .in(wire_28), .out(wire_70_26));
  TC_Switch # (.UUID(64'd1920741343055373206 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_353 (.en(wire_209), .in(wire_37), .out(wire_70_27));
  TC_Switch # (.UUID(64'd4021669768454360472 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_354 (.en(wire_65), .in(wire_96), .out(wire_70_28));
  TC_Switch # (.UUID(64'd1889670277106741446 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_355 (.en(wire_160), .in(wire_3), .out(wire_70_29));
  TC_Switch # (.UUID(64'd3260985352587339952 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_356 (.en(wire_425), .in(wire_150), .out(wire_70_30));
  TC_Switch # (.UUID(64'd2575338778244414098 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_357 (.en(wire_272), .in(wire_221), .out(wire_70_31));
  TC_Splitter8 # (.UUID(64'd4330732377258575308 ^ UUID)) Splitter8_358 (.in(wire_199), .out0(wire_188), .out1(wire_11), .out2(wire_122), .out3(wire_209), .out4(wire_65), .out5(wire_160), .out6(wire_425), .out7(wire_272));
  TC_Buffer # (.UUID(64'd203309114433716697 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_359 (.in(wire_167), .out(wire_15));
  TC_Buffer # (.UUID(64'd4497935948046771375 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_360 (.in(wire_70), .out(wire_256));
  TC_Constant # (.UUID(64'd2652289593323316064 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h0)) Constant32_361 (.out(wire_311));
  TC_Buffer # (.UUID(64'd3403365156378003067 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_362 (.in(wire_107), .out(wire_355));
  TC_Buffer # (.UUID(64'd2078592390335996446 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_363 (.in(wire_1), .out());
  TC_Buffer # (.UUID(64'd779922314171047114 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_364 (.in(wire_53), .out(wire_409));
  TC_Buffer # (.UUID(64'd149917869844955214 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_365 (.in(wire_214), .out(wire_313));
  TC_Buffer # (.UUID(64'd3148727733132701959 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_366 (.in(wire_176), .out(wire_385));
  TC_Buffer # (.UUID(64'd4478883126463910117 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_367 (.in(wire_135), .out(wire_131));
  TC_Buffer # (.UUID(64'd1509087869747369071 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_368 (.in(wire_118), .out(wire_339));
  TC_Buffer # (.UUID(64'd3078292029986845944 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_369 (.in(wire_173), .out(wire_285));
  TC_Buffer # (.UUID(64'd2931833856900649059 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_370 (.in(wire_45), .out(wire_191));
  TC_Buffer # (.UUID(64'd3580487990483905896 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_371 (.in(wire_215), .out(wire_421));
  TC_Buffer # (.UUID(64'd1147538542811540042 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_372 (.in(wire_162), .out(wire_408));
  TC_Buffer # (.UUID(64'd826894211383350680 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_373 (.in(wire_116), .out(wire_284));
  TC_Buffer # (.UUID(64'd3771532439236542689 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_374 (.in(wire_126), .out(wire_60));
  TC_Buffer # (.UUID(64'd853044613490682130 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_375 (.in(wire_198), .out(wire_353));
  TC_Buffer # (.UUID(64'd1230146387499610852 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_376 (.in(wire_88), .out(wire_17));
  TC_Buffer # (.UUID(64'd1156530599392149419 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_377 (.in(wire_228), .out(wire_18));
  TC_Buffer # (.UUID(64'd1385870454688759788 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_378 (.in(wire_111), .out(wire_379));
  TC_Buffer # (.UUID(64'd435724858089039808 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_379 (.in(wire_99), .out(wire_386));
  TC_Buffer # (.UUID(64'd2358704279662367987 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_380 (.in(wire_63), .out(wire_336));
  TC_Buffer # (.UUID(64'd473881130067592486 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_381 (.in(wire_267), .out(wire_211));
  TC_Buffer # (.UUID(64'd341597032268246022 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_382 (.in(wire_95), .out(wire_444));
  TC_Buffer # (.UUID(64'd722725231027671654 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_383 (.in(wire_179), .out(wire_246));
  TC_Buffer # (.UUID(64'd4475455387665777511 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_384 (.in(wire_21), .out(wire_113));
  TC_Buffer # (.UUID(64'd809532325430816339 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_385 (.in(wire_128), .out(wire_330));
  TC_Buffer # (.UUID(64'd3225970828693863241 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_386 (.in(wire_159), .out(wire_365));
  TC_Buffer # (.UUID(64'd1713264642969941712 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_387 (.in(wire_110), .out(wire_233));
  TC_Buffer # (.UUID(64'd246997092383671131 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_388 (.in(wire_249), .out(wire_264));
  TC_Buffer # (.UUID(64'd3561534574736112586 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_389 (.in(wire_28), .out(wire_295));
  TC_Buffer # (.UUID(64'd349573961585296007 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_390 (.in(wire_37), .out(wire_251));
  TC_Buffer # (.UUID(64'd1370175540667521266 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_391 (.in(wire_96), .out(wire_181));
  TC_Buffer # (.UUID(64'd4577111249699879360 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_392 (.in(wire_3), .out(wire_376));
  TC_Buffer # (.UUID(64'd2445382406320351400 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_393 (.in(wire_150), .out(wire_297));
  TC_Buffer # (.UUID(64'd781538958166454725 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_394 (.in(wire_221), .out(wire_125));
  TC_Maker8 # (.UUID(64'd3488007923077716303 ^ UUID)) Maker8_395 (.in0(wire_288), .in1(wire_340), .in2(wire_102), .in3(wire_195), .in4(wire_71), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_117));
  TC_Maker8 # (.UUID(64'd1833178259065145121 ^ UUID)) Maker8_396 (.in0(wire_84), .in1(wire_332), .in2(wire_220), .in3(wire_301), .in4(wire_449), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_203));
  TC_Maker8 # (.UUID(64'd4057909194347133542 ^ UUID)) Maker8_397 (.in0(wire_364), .in1(wire_382), .in2(wire_158), .in3(wire_343), .in4(wire_363), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_155));
  TC_Constant # (.UUID(64'd1266887650110149333 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_398 (.out(wire_87));
  TC_Shl # (.UUID(64'd3860679339152863391 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_399 (.in({{31{1'b0}}, wire_87 }), .shift(wire_117), .out(wire_78));
  TC_Constant # (.UUID(64'd3110180527670241762 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_400 (.out(wire_438));
  TC_Shl # (.UUID(64'd3770848241066039869 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_401 (.in({{31{1'b0}}, wire_438 }), .shift(wire_203), .out(wire_315));
  TC_Constant # (.UUID(64'd2101249925536989277 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_402 (.out(wire_342));
  TC_Shl # (.UUID(64'd1748919223126118636 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_403 (.in({{31{1'b0}}, wire_342 }), .shift(wire_155), .out(wire_432));
  TC_Buffer # (.UUID(64'd2824446733315679492 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_404 (.in(wire_115), .out(wire_351));
  TC_Buffer # (.UUID(64'd3742829896238883482 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_405 (.in(wire_231), .out(wire_362));
  TC_Buffer # (.UUID(64'd2724346673473456697 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_406 (.in(wire_9), .out(wire_255));
  TC_Buffer # (.UUID(64'd4429420174311818155 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_407 (.in(wire_62), .out(wire_208));
  TC_Buffer # (.UUID(64'd3161096343730813467 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_408 (.in(wire_427), .out(wire_25));
  TC_Buffer # (.UUID(64'd4080693366154061052 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_409 (.in(wire_73), .out(wire_241));
  TC_Shr # (.UUID(64'd768819421975172603 ^ UUID), .BIT_WIDTH(64'd64)) Shr64_410 (.in(wire_208), .shift(wire_422), .out(wire_427));
  TC_Constant # (.UUID(64'd2185369399685244588 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_411 (.out(wire_422));
  TC_And # (.UUID(64'd1674364192246079449 ^ UUID), .BIT_WIDTH(64'd64)) And64_412 (.in0(wire_208), .in1(wire_156), .out(wire_269));
  TC_Constant # (.UUID(64'd3213227198313095996 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h7)) Constant64_413 (.out(wire_156));
  TC_Buffer # (.UUID(64'd925811751658486003 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_414 (.in(wire_154), .out(wire_109));
  TC_Shr # (.UUID(64'd1364216107044831048 ^ UUID), .BIT_WIDTH(64'd64)) Shr64_415 (.in(wire_280), .shift(wire_81), .out(wire_154));
  TC_And # (.UUID(64'd2639533957149927325 ^ UUID), .BIT_WIDTH(64'd64)) And64_416 (.in0(wire_29), .in1(wire_388), .out(wire_280));
  TC_Not # (.UUID(64'd2391628148256969402 ^ UUID), .BIT_WIDTH(64'd64)) Not64_417 (.in(wire_324), .out(wire_424));
  TC_And # (.UUID(64'd122266305254588552 ^ UUID), .BIT_WIDTH(64'd64)) And64_418 (.in0(wire_424), .in1(wire_29), .out(wire_394));
  TC_Or # (.UUID(64'd237919812159994493 ^ UUID), .BIT_WIDTH(64'd64)) Or64_419 (.in0(wire_43), .in1(wire_394), .out(wire_73));
  TC_And # (.UUID(64'd1717030403840026689 ^ UUID), .BIT_WIDTH(64'd64)) And64_420 (.in0(wire_255), .in1(wire_193), .out(wire_419));
  TC_Buffer # (.UUID(64'd187451873155405380 ^ UUID), .BIT_WIDTH(64'd64)) Buffer64_421 (.in(wire_29), .out());
  TC_Shl # (.UUID(64'd2257392532296178393 ^ UUID), .BIT_WIDTH(64'd64)) Shl64_422 (.in(wire_273), .shift(wire_81), .out(wire_388));
  TC_Shl # (.UUID(64'd3452680584397757071 ^ UUID), .BIT_WIDTH(64'd64)) Shl64_423 (.in(wire_193), .shift(wire_81), .out(wire_324));
  TC_Shl # (.UUID(64'd562267020645338885 ^ UUID), .BIT_WIDTH(64'd64)) Shl64_424 (.in(wire_419), .shift(wire_81), .out(wire_43));
  _64bitz_Selector # (.UUID(64'd837285822481470997 ^ UUID)) _64bitz_Selector_425 (.clk(clk), .rst(rst), .Bytes(wire_362), .Output(wire_273));
  _64bitz_Selector # (.UUID(64'd3236062019093102112 ^ UUID)) _64bitz_Selector_426 (.clk(clk), .rst(rst), .Bytes(wire_351), .Output(wire_193));
  TC_Shl # (.UUID(64'd263565130673154455 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_427 (.in(wire_269[7:0]), .shift(wire_439), .out(wire_81));
  TC_Constant # (.UUID(64'd43642452680328666 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_428 (.out(wire_439));
  TC_Buffer # (.UUID(64'd3442681514873585622 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_429 (.in(wire_15), .out(wire_145));
  TC_Buffer # (.UUID(64'd814663592506655634 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_430 (.in(wire_256), .out(wire_48));
  TC_Buffer # (.UUID(64'd4192911053225322289 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_431 (.in(wire_141), .out(wire_258));
  TC_Switch # (.UUID(64'd3008015254934111552 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_432 (.en(wire_367), .in(wire_123), .out(wire_1_2));
  TC_Splitter32 # (.UUID(64'd1450832447418184470 ^ UUID)) Splitter32_433 (.in(wire_168), .out0(wire_435), .out1(wire_180), .out2(), .out3());
  TC_Splitter8 # (.UUID(64'd569486895244707668 ^ UUID)) Splitter8_434 (.in(wire_435), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(wire_130), .out6(), .out7());
  TC_Buffer # (.UUID(64'd121554546992970759 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_435 (.in(wire_105), .out(wire_142));
  TC_Splitter8 # (.UUID(64'd442772438262865453 ^ UUID)) Splitter8_436 (.in(wire_180), .out0(), .out1(), .out2(), .out3(), .out4(wire_279), .out5(wire_67), .out6(wire_114), .out7());
  TC_Decoder3 # (.UUID(64'd2173384068657890044 ^ UUID)) Decoder3_437 (.dis(1'd0), .sel0(wire_279), .sel1(wire_67), .sel2(wire_114), .out0(wire_146), .out1(wire_348), .out2(wire_31), .out3(wire_6), .out4(wire_245), .out5(wire_121), .out6(wire_434), .out7(wire_119));
  TC_Ashr # (.UUID(64'd4519441965371985183 ^ UUID), .BIT_WIDTH(64'd32)) Ashr32_438 (.in(wire_168), .shift(wire_291), .out(wire_186));
  TC_Constant # (.UUID(64'd2553359768039302569 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h14)) Constant8_439 (.out(wire_291));
  TC_Ashr # (.UUID(64'd1938985463505896238 ^ UUID), .BIT_WIDTH(64'd32)) Ashr32_440 (.in(wire_168), .shift(wire_445), .out(wire_305));
  TC_Constant # (.UUID(64'd2113505211085757844 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h19)) Constant8_441 (.out(wire_445));
  TC_Add # (.UUID(64'd1806826801169682507 ^ UUID), .BIT_WIDTH(64'd32)) Add32_442 (.in0(wire_145), .in1(wire_186), .ci(1'd0), .out(wire_350), .co());
  TC_Buffer # (.UUID(64'd3296931108182422958 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_443 (.in(wire_429[7:0]), .out(wire_306));
  TC_Switch # (.UUID(64'd3188424604856445666 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_444 (.en(wire_146), .in(wire_359), .out(wire_169_3));
  TC_Splitter32 # (.UUID(64'd4298750993472201539 ^ UUID)) Splitter32_445 (.in(wire_19), .out0(wire_372), .out1(), .out2(), .out3());
  TC_Splitter8 # (.UUID(64'd1132354071000996356 ^ UUID)) Splitter8_446 (.in(wire_372), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_13));
  TC_Maker32 # (.UUID(64'd1893638985581802478 ^ UUID)) Maker32_447 (.in0(wire_372), .in1(wire_172), .in2(wire_172), .in3(wire_172), .out(wire_359));
  TC_Maker8 # (.UUID(64'd2505817213189423649 ^ UUID)) Maker8_448 (.in0(wire_13), .in1(wire_13), .in2(wire_13), .in3(wire_13), .in4(wire_13), .in5(wire_13), .in6(wire_13), .in7(wire_13), .out(wire_172));
  TC_Splitter32 # (.UUID(64'd4103965242347969359 ^ UUID)) Splitter32_449 (.in(wire_19), .out0(wire_254), .out1(wire_40), .out2(), .out3());
  TC_Splitter8 # (.UUID(64'd2083671351688561564 ^ UUID)) Splitter8_450 (.in(wire_40), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_4));
  TC_Maker8 # (.UUID(64'd1795792930892414866 ^ UUID)) Maker8_451 (.in0(wire_4), .in1(wire_4), .in2(wire_4), .in3(wire_4), .in4(wire_4), .in5(wire_4), .in6(wire_4), .in7(wire_4), .out(wire_300));
  TC_Maker32 # (.UUID(64'd206357386023687990 ^ UUID)) Maker32_452 (.in0(wire_254), .in1(wire_40), .in2(wire_300), .in3(wire_300), .out(wire_393));
  TC_Switch # (.UUID(64'd2283289723681929728 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_453 (.en(wire_348), .in(wire_393), .out(wire_169_0));
  TC_Switch # (.UUID(64'd1578447547286228622 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_454 (.en(wire_31), .in(wire_19), .out(wire_169_1));
  TC_Switch # (.UUID(64'd3791668145762299402 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_455 (.en(wire_245), .in(wire_378), .out(wire_169_2));
  TC_Switch # (.UUID(64'd4554041588454622461 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_456 (.en(wire_121), .in(wire_8), .out(wire_169_4));
  TC_Add # (.UUID(64'd1625149425280856650 ^ UUID), .BIT_WIDTH(64'd32)) Add32_457 (.in0(wire_145), .in1(wire_260), .ci(1'd0), .out(wire_20), .co());
  TC_Shl # (.UUID(64'd3282922818602697939 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_458 (.in(wire_305), .shift(wire_443), .out(wire_304));
  TC_Constant # (.UUID(64'd3942845999438537981 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_459 (.out(wire_443));
  TC_Or # (.UUID(64'd2735627082527286231 ^ UUID), .BIT_WIDTH(64'd32)) Or32_460 (.in0(wire_304), .in1(wire_265), .out(wire_260));
  TC_Shr # (.UUID(64'd839122501473322725 ^ UUID), .BIT_WIDTH(64'd32)) Shr32_461 (.in(wire_168), .shift(wire_433), .out(wire_75));
  TC_Constant # (.UUID(64'd3308612162966646265 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_462 (.out(wire_433));
  TC_Constant # (.UUID(64'd2823609753204562993 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_463 (.out(wire_399));
  TC_And # (.UUID(64'd2617873379414410143 ^ UUID), .BIT_WIDTH(64'd32)) And32_464 (.in0(wire_75), .in1({{24{1'b0}}, wire_399 }), .out(wire_265));
  TC_Decoder3 # (.UUID(64'd350899084139630687 ^ UUID)) Decoder3_465 (.dis(1'd0), .sel0(wire_279), .sel1(wire_67), .sel2(wire_114), .out0(wire_171), .out1(wire_328), .out2(wire_222), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd1812732707729274731 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_466 (.en(wire_171), .in(wire_392), .out(wire_247_0));
  TC_Constant # (.UUID(64'd3738910968182952104 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_467 (.out(wire_392));
  TC_Switch # (.UUID(64'd4067772386914195036 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_468 (.en(wire_328), .in(wire_190), .out(wire_247_1));
  TC_Constant # (.UUID(64'd1605021603375967928 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_469 (.out(wire_190));
  TC_Switch # (.UUID(64'd1730122275101123611 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_470 (.en(wire_222), .in(wire_371), .out(wire_247_2));
  TC_Constant # (.UUID(64'd1715468856498864266 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_471 (.out(wire_371));
  TC_Constant # (.UUID(64'd2976333720201650127 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_472 (.out(wire_192));
  TC_Switch # (.UUID(64'd2209381333052485081 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_473 (.en(wire_366), .in(wire_192), .out(wire_184_0));
  TC_Or # (.UUID(64'd1994103989963715350 ^ UUID), .BIT_WIDTH(64'd1)) Or_474 (.in0(wire_146), .in1(wire_245), .out(wire_366));
  TC_Constant # (.UUID(64'd1358490902349266189 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_475 (.out(wire_144));
  TC_Switch # (.UUID(64'd4299599623468776896 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_476 (.en(wire_441), .in(wire_144), .out(wire_184_1));
  TC_Or # (.UUID(64'd4012036525874190182 ^ UUID), .BIT_WIDTH(64'd1)) Or_477 (.in0(wire_348), .in1(wire_121), .out(wire_441));
  TC_Constant # (.UUID(64'd2358578198838993326 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_478 (.out(wire_396));
  TC_Switch # (.UUID(64'd1025812563839059013 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_479 (.en(wire_31), .in(wire_396), .out(wire_184_2));
  TC_Not # (.UUID(64'd1954730347310721103 ^ UUID), .BIT_WIDTH(64'd1)) Not_480 (.in(wire_130), .out(wire_296));
  TC_Constant # (.UUID(64'd3989431052611746113 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_481 (.out(wire_187));
  TC_Switch # (.UUID(64'd1419455945234160340 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_482 (.en(wire_258), .in(wire_296), .out(wire_56));
  TC_Switch # (.UUID(64'd1182382243167072162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_483 (.en(wire_258), .in(wire_130), .out(wire_257));
  TC_DelayLine # (.UUID(64'd868337229697359879 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_484 (.clk(clk), .rst(rst), .in(wire_257), .out(wire_7));
  TC_DelayLine # (.UUID(64'd3074871992927228768 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_485 (.clk(clk), .rst(rst), .in(wire_56), .out(wire_143));
  TC_Buffer # (.UUID(64'd3076301426948079881 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_486 (.in(wire_143), .out(wire_314));
  TC_Mux # (.UUID(64'd3294096435622679339 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_487 (.sel(wire_7), .in0(wire_169), .in1(wire_48), .out(wire_123));
  TC_Or # (.UUID(64'd1874480084249769784 ^ UUID), .BIT_WIDTH(64'd1)) Or_488 (.in0(wire_7), .in1(wire_143), .out(wire_367));
  TC_Nor # (.UUID(64'd275282978308376820 ^ UUID), .BIT_WIDTH(64'd1)) Nor_489 (.in0(wire_7), .in1(wire_143), .out(wire_283));
  TC_DelayLine # (.UUID(64'd88320780327091975 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_490 (.clk(clk), .rst(rst), .in(wire_168), .out(wire_147));
  TC_Mux # (.UUID(64'd2285835871575853886 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_491 (.sel(wire_242), .in0(wire_184), .in1(wire_187), .out(wire_69));
  TC_Buffer # (.UUID(64'd2068176701917864040 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_492 (.in(wire_147), .out(wire_174));
  TC_Switch # (.UUID(64'd3398197759057014925 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_493 (.en(wire_7), .in({{24{1'b0}}, wire_247 }), .out(wire_429));
  TC_Buffer # (.UUID(64'd4117688863481788720 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_494 (.in(wire_333), .out(wire_108));
  TC_Not # (.UUID(64'd348338904957669946 ^ UUID), .BIT_WIDTH(64'd1)) Not_495 (.in(wire_56), .out(wire_242));
  TC_DelayLine # (.UUID(64'd72091540950518397 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_496 (.clk(clk), .rst(rst), .in(wire_69), .out(wire_333));
  TC_Buffer # (.UUID(64'd1258988992638853442 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_497 (.in(wire_283), .out(wire_182));
  TC_Buffer # (.UUID(64'd2001413141544554488 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_498 (.in(wire_243), .out(wire_168));
  TC_DelayLine # (.UUID(64'd2881589807745929050 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_499 (.clk(clk), .rst(rst), .in(wire_350), .out(wire_129));
  TC_DelayLine # (.UUID(64'd597166326161706409 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_500 (.clk(clk), .rst(rst), .in(wire_20), .out(wire_46));
  TC_Buffer # (.UUID(64'd4156479662433209742 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_501 (.in(wire_436), .out(wire_33));
  TC_Buffer # (.UUID(64'd2418485793995780281 ^ UUID), .BIT_WIDTH(64'd32)) Buffer32_502 (.in(wire_109[31:0]), .out(wire_19));
  TC_Constant # (.UUID(64'd322763907399541861 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFF)) Constant32_503 (.out(wire_344));
  TC_Constant # (.UUID(64'd3235559750950740763 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFFFF)) Constant32_504 (.out(wire_430));
  TC_And # (.UUID(64'd3520851976516274068 ^ UUID), .BIT_WIDTH(64'd32)) And32_505 (.in0(wire_19), .in1(wire_344), .out(wire_378));
  TC_And # (.UUID(64'd2130438836809759628 ^ UUID), .BIT_WIDTH(64'd32)) And32_506 (.in0(wire_19), .in1(wire_430), .out(wire_8));
  TC_Or # (.UUID(64'd4523391179892267281 ^ UUID), .BIT_WIDTH(64'd1)) Or_507 (.in0(wire_7), .in1(wire_143), .out(wire_389));
  _2z_Wayz_Switch # (.UUID(64'd2532554746192223676 ^ UUID)) _2z_Wayz_Switch_508 (.clk(clk), .rst(rst), .Input_1(wire_143), .Input_2(wire_7), .Input_3(wire_142), .Input_4(wire_46), .Input_5(wire_129), .Input_6(32'd0), .Output(wire_436));

  wire [63:0] wire_0;
  wire [31:0] wire_1;
  wire [31:0] wire_1_0;
  wire [31:0] wire_1_1;
  wire [31:0] wire_1_2;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2;
  wire [63:0] wire_2;
  wire [31:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [31:0] wire_8;
  wire [63:0] wire_9;
  wire [31:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [31:0] wire_14;
  wire [31:0] wire_15;
  wire [0:0] wire_16;
  wire [31:0] wire_17;
  wire [31:0] wire_18;
  wire [31:0] wire_19;
  wire [31:0] wire_20;
  wire [31:0] wire_21;
  wire [31:0] wire_22;
  wire [31:0] wire_23;
  wire [63:0] wire_24;
  wire [63:0] wire_25;
  wire [63:0] wire_26;
  wire [0:0] wire_27;
  wire [31:0] wire_28;
  wire [63:0] wire_29;
  wire [63:0] wire_29_0;
  wire [63:0] wire_29_1;
  wire [63:0] wire_29_2;
  assign wire_29 = wire_29_0|wire_29_1|wire_29_2;
  wire [63:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [31:0] wire_33;
  wire [31:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [31:0] wire_37;
  wire [31:0] wire_38;
  wire [31:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [63:0] wire_42;
  wire [63:0] wire_43;
  wire [63:0] wire_44;
  wire [31:0] wire_45;
  wire [31:0] wire_46;
  wire [0:0] wire_47;
  wire [31:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [31:0] wire_52;
  wire [31:0] wire_53;
  wire [0:0] wire_54;
  wire [31:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [31:0] wire_58;
  wire [0:0] wire_59;
  wire [31:0] wire_60;
  wire [0:0] wire_61;
  wire [63:0] wire_62;
  wire [31:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [63:0] wire_66;
  wire [0:0] wire_67;
  wire [31:0] wire_68;
  wire [7:0] wire_69;
  wire [31:0] wire_70;
  wire [31:0] wire_70_0;
  wire [31:0] wire_70_1;
  wire [31:0] wire_70_2;
  wire [31:0] wire_70_3;
  wire [31:0] wire_70_4;
  wire [31:0] wire_70_5;
  wire [31:0] wire_70_6;
  wire [31:0] wire_70_7;
  wire [31:0] wire_70_8;
  wire [31:0] wire_70_9;
  wire [31:0] wire_70_10;
  wire [31:0] wire_70_11;
  wire [31:0] wire_70_12;
  wire [31:0] wire_70_13;
  wire [31:0] wire_70_14;
  wire [31:0] wire_70_15;
  wire [31:0] wire_70_16;
  wire [31:0] wire_70_17;
  wire [31:0] wire_70_18;
  wire [31:0] wire_70_19;
  wire [31:0] wire_70_20;
  wire [31:0] wire_70_21;
  wire [31:0] wire_70_22;
  wire [31:0] wire_70_23;
  wire [31:0] wire_70_24;
  wire [31:0] wire_70_25;
  wire [31:0] wire_70_26;
  wire [31:0] wire_70_27;
  wire [31:0] wire_70_28;
  wire [31:0] wire_70_29;
  wire [31:0] wire_70_30;
  wire [31:0] wire_70_31;
  assign wire_70 = wire_70_0|wire_70_1|wire_70_2|wire_70_3|wire_70_4|wire_70_5|wire_70_6|wire_70_7|wire_70_8|wire_70_9|wire_70_10|wire_70_11|wire_70_12|wire_70_13|wire_70_14|wire_70_15|wire_70_16|wire_70_17|wire_70_18|wire_70_19|wire_70_20|wire_70_21|wire_70_22|wire_70_23|wire_70_24|wire_70_25|wire_70_26|wire_70_27|wire_70_28|wire_70_29|wire_70_30|wire_70_31;
  wire [0:0] wire_71;
  wire [7:0] wire_72;
  wire [63:0] wire_73;
  wire [7:0] wire_74;
  wire [31:0] wire_75;
  wire [31:0] wire_76;
  wire [0:0] wire_77;
  wire [31:0] wire_78;
  wire [31:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [7:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [31:0] wire_85;
  wire [31:0] wire_86;
  wire [0:0] wire_87;
  wire [31:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [63:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [31:0] wire_95;
  wire [31:0] wire_96;
  wire [0:0] wire_97;
  wire [63:0] wire_98;
  wire [31:0] wire_99;
  wire [63:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [63:0] wire_104;
  wire [31:0] wire_105;
  wire [31:0] wire_106;
  wire [0:0] wire_107;
  wire [7:0] wire_108;
  wire [63:0] wire_109;
  wire [31:0] wire_110;
  wire [31:0] wire_111;
  wire [0:0] wire_112;
  wire [31:0] wire_113;
  wire [0:0] wire_114;
  wire [7:0] wire_115;
  wire [31:0] wire_116;
  wire [7:0] wire_117;
  wire [31:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [31:0] wire_123;
  wire [0:0] wire_124;
  wire [31:0] wire_125;
  wire [31:0] wire_126;
  wire [0:0] wire_127;
  wire [31:0] wire_128;
  wire [31:0] wire_129;
  wire [0:0] wire_130;
  wire [31:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [31:0] wire_135;
  wire [63:0] wire_136;
  wire [31:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [0:0] wire_141;
  wire [31:0] wire_142;
  wire [0:0] wire_143;
  wire [7:0] wire_144;
  wire [31:0] wire_145;
  wire [0:0] wire_146;
  wire [31:0] wire_147;
  wire [7:0] wire_148;
  wire [0:0] wire_149;
  wire [31:0] wire_150;
  wire [0:0] wire_151;
  wire [0:0] wire_152;
  wire [0:0] wire_153;
  wire [63:0] wire_154;
  wire [7:0] wire_155;
  wire [63:0] wire_156;
  wire [0:0] wire_157;
  wire [0:0] wire_158;
  wire [31:0] wire_159;
  wire [0:0] wire_160;
  wire [0:0] wire_161;
  wire [31:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [0:0] wire_165;
  wire [0:0] wire_166;
  wire [31:0] wire_167;
  wire [31:0] wire_167_0;
  wire [31:0] wire_167_1;
  wire [31:0] wire_167_2;
  wire [31:0] wire_167_3;
  wire [31:0] wire_167_4;
  wire [31:0] wire_167_5;
  wire [31:0] wire_167_6;
  wire [31:0] wire_167_7;
  wire [31:0] wire_167_8;
  wire [31:0] wire_167_9;
  wire [31:0] wire_167_10;
  wire [31:0] wire_167_11;
  wire [31:0] wire_167_12;
  wire [31:0] wire_167_13;
  wire [31:0] wire_167_14;
  wire [31:0] wire_167_15;
  wire [31:0] wire_167_16;
  wire [31:0] wire_167_17;
  wire [31:0] wire_167_18;
  wire [31:0] wire_167_19;
  wire [31:0] wire_167_20;
  wire [31:0] wire_167_21;
  wire [31:0] wire_167_22;
  wire [31:0] wire_167_23;
  wire [31:0] wire_167_24;
  wire [31:0] wire_167_25;
  wire [31:0] wire_167_26;
  wire [31:0] wire_167_27;
  wire [31:0] wire_167_28;
  wire [31:0] wire_167_29;
  wire [31:0] wire_167_30;
  wire [31:0] wire_167_31;
  assign wire_167 = wire_167_0|wire_167_1|wire_167_2|wire_167_3|wire_167_4|wire_167_5|wire_167_6|wire_167_7|wire_167_8|wire_167_9|wire_167_10|wire_167_11|wire_167_12|wire_167_13|wire_167_14|wire_167_15|wire_167_16|wire_167_17|wire_167_18|wire_167_19|wire_167_20|wire_167_21|wire_167_22|wire_167_23|wire_167_24|wire_167_25|wire_167_26|wire_167_27|wire_167_28|wire_167_29|wire_167_30|wire_167_31;
  wire [31:0] wire_168;
  wire [31:0] wire_169;
  wire [31:0] wire_169_0;
  wire [31:0] wire_169_1;
  wire [31:0] wire_169_2;
  wire [31:0] wire_169_3;
  wire [31:0] wire_169_4;
  assign wire_169 = wire_169_0|wire_169_1|wire_169_2|wire_169_3|wire_169_4;
  wire [0:0] wire_170;
  wire [0:0] wire_171;
  wire [7:0] wire_172;
  wire [31:0] wire_173;
  wire [31:0] wire_174;
  wire [0:0] wire_175;
  wire [31:0] wire_176;
  wire [0:0] wire_177;
  wire [0:0] wire_178;
  wire [31:0] wire_179;
  wire [7:0] wire_180;
  wire [31:0] wire_181;
  wire [0:0] wire_182;
  wire [0:0] wire_183;
  wire [7:0] wire_184;
  wire [7:0] wire_184_0;
  wire [7:0] wire_184_1;
  wire [7:0] wire_184_2;
  assign wire_184 = wire_184_0|wire_184_1|wire_184_2;
  wire [0:0] wire_185;
  wire [31:0] wire_186;
  wire [7:0] wire_187;
  wire [0:0] wire_188;
  wire [0:0] wire_189;
  wire [7:0] wire_190;
  wire [31:0] wire_191;
  wire [7:0] wire_192;
  wire [63:0] wire_193;
  wire [0:0] wire_194;
  wire [0:0] wire_195;
  wire [0:0] wire_196;
  wire [0:0] wire_197;
  wire [31:0] wire_198;
  wire [7:0] wire_199;
  wire [0:0] wire_200;
  wire [7:0] wire_201;
  wire [0:0] wire_202;
  wire [7:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [0:0] wire_206;
  wire [0:0] wire_207;
  wire [63:0] wire_208;
  wire [0:0] wire_209;
  wire [0:0] wire_210;
  wire [31:0] wire_211;
  wire [0:0] wire_212;
  wire [7:0] wire_213;
  wire [31:0] wire_214;
  wire [31:0] wire_215;
  wire [7:0] wire_216;
  wire [7:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [31:0] wire_221;
  wire [0:0] wire_222;
  wire [0:0] wire_223;
  wire [7:0] wire_224;
  wire [0:0] wire_225;
  wire [0:0] wire_226;
  wire [31:0] wire_227;
  wire [31:0] wire_228;
  wire [0:0] wire_229;
  wire [0:0] wire_230;
  wire [7:0] wire_231;
  wire [63:0] wire_232;
  wire [31:0] wire_233;
  wire [0:0] wire_234;
  wire [0:0] wire_235;
  wire [0:0] wire_236;
  wire [0:0] wire_237;
  wire [0:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [63:0] wire_241;
  wire [0:0] wire_242;
  wire [31:0] wire_243;
  wire [0:0] wire_244;
  wire [0:0] wire_245;
  wire [31:0] wire_246;
  wire [7:0] wire_247;
  wire [7:0] wire_247_0;
  wire [7:0] wire_247_1;
  wire [7:0] wire_247_2;
  assign wire_247 = wire_247_0|wire_247_1|wire_247_2;
  wire [0:0] wire_248;
  wire [31:0] wire_249;
  wire [0:0] wire_250;
  wire [31:0] wire_251;
  wire [0:0] wire_252;
  wire [0:0] wire_253;
  wire [7:0] wire_254;
  wire [63:0] wire_255;
  wire [31:0] wire_256;
  wire [0:0] wire_257;
  wire [0:0] wire_258;
  wire [0:0] wire_259;
  wire [31:0] wire_260;
  wire [0:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [31:0] wire_264;
  wire [31:0] wire_265;
  wire [0:0] wire_266;
  wire [31:0] wire_267;
  wire [0:0] wire_268;
  assign wire_268 = 0;
  wire [63:0] wire_269;
  wire [0:0] wire_270;
  wire [0:0] wire_271;
  wire [0:0] wire_272;
  wire [63:0] wire_273;
  wire [7:0] wire_274;
  wire [7:0] wire_275;
  wire [0:0] wire_276;
  wire [7:0] wire_277;
  wire [0:0] wire_278;
  wire [0:0] wire_279;
  wire [63:0] wire_280;
  wire [0:0] wire_281;
  wire [0:0] wire_282;
  wire [0:0] wire_283;
  wire [31:0] wire_284;
  wire [31:0] wire_285;
  wire [0:0] wire_286;
  wire [0:0] wire_287;
  wire [0:0] wire_288;
  wire [0:0] wire_289;
  wire [0:0] wire_290;
  wire [7:0] wire_291;
  wire [0:0] wire_292;
  wire [31:0] wire_293;
  wire [0:0] wire_294;
  wire [31:0] wire_295;
  wire [0:0] wire_296;
  wire [31:0] wire_297;
  wire [7:0] wire_298;
  wire [0:0] wire_299;
  wire [7:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [0:0] wire_303;
  wire [31:0] wire_304;
  wire [31:0] wire_305;
  wire [7:0] wire_306;
  wire [0:0] wire_307;
  wire [0:0] wire_308;
  wire [0:0] wire_309;
  wire [63:0] wire_310;
  wire [31:0] wire_311;
  wire [0:0] wire_312;
  wire [31:0] wire_313;
  wire [0:0] wire_314;
  wire [31:0] wire_315;
  wire [7:0] wire_316;
  wire [0:0] wire_317;
  wire [7:0] wire_318;
  wire [7:0] wire_319;
  wire [0:0] wire_320;
  wire [7:0] wire_321;
  wire [31:0] wire_322;
  wire [63:0] wire_323;
  wire [63:0] wire_324;
  wire [31:0] wire_325;
  wire [7:0] wire_326;
  wire [0:0] wire_327;
  wire [0:0] wire_328;
  wire [31:0] wire_329;
  wire [31:0] wire_330;
  wire [7:0] wire_331;
  wire [0:0] wire_332;
  wire [7:0] wire_333;
  wire [0:0] wire_334;
  wire [0:0] wire_335;
  wire [31:0] wire_336;
  wire [0:0] wire_337;
  assign wire_337 = 0;
  wire [63:0] wire_338;
  wire [31:0] wire_339;
  wire [0:0] wire_340;
  wire [0:0] wire_341;
  assign wire_341 = 0;
  wire [0:0] wire_342;
  wire [0:0] wire_343;
  wire [31:0] wire_344;
  wire [63:0] wire_345;
  wire [63:0] wire_346;
  wire [0:0] wire_347;
  wire [0:0] wire_348;
  wire [0:0] wire_349;
  wire [31:0] wire_350;
  wire [7:0] wire_351;
  wire [0:0] wire_352;
  wire [31:0] wire_353;
  wire [0:0] wire_354;
  wire [0:0] wire_355;
  wire [0:0] wire_356;
  wire [0:0] wire_357;
  wire [0:0] wire_358;
  wire [31:0] wire_359;
  wire [0:0] wire_360;
  wire [0:0] wire_361;
  wire [7:0] wire_362;
  wire [0:0] wire_363;
  wire [0:0] wire_364;
  wire [31:0] wire_365;
  wire [0:0] wire_366;
  wire [0:0] wire_367;
  wire [0:0] wire_368;
  wire [15:0] wire_369;
  wire [0:0] wire_370;
  wire [7:0] wire_371;
  wire [7:0] wire_372;
  wire [0:0] wire_373;
  wire [0:0] wire_374;
  wire [0:0] wire_375;
  wire [31:0] wire_376;
  wire [0:0] wire_377;
  wire [31:0] wire_378;
  wire [31:0] wire_379;
  wire [0:0] wire_380;
  wire [0:0] wire_381;
  wire [0:0] wire_382;
  wire [63:0] wire_383;
  wire [0:0] wire_384;
  wire [31:0] wire_385;
  wire [31:0] wire_386;
  wire [0:0] wire_387;
  wire [63:0] wire_388;
  wire [0:0] wire_389;
  wire [0:0] wire_390;
  wire [0:0] wire_391;
  wire [7:0] wire_392;
  wire [31:0] wire_393;
  wire [63:0] wire_394;
  wire [0:0] wire_395;
  wire [7:0] wire_396;
  wire [0:0] wire_397;
  wire [0:0] wire_398;
  wire [7:0] wire_399;
  wire [63:0] wire_400;
  wire [0:0] wire_401;
  wire [0:0] wire_402;
  wire [0:0] wire_403;
  wire [0:0] wire_404;
  wire [0:0] wire_405;
  wire [0:0] wire_406;
  wire [0:0] wire_407;
  wire [31:0] wire_408;
  wire [31:0] wire_409;
  wire [0:0] wire_410;
  wire [63:0] wire_411;
  wire [0:0] wire_412;
  wire [0:0] wire_413;
  wire [63:0] wire_414;
  wire [7:0] wire_415;
  wire [63:0] wire_416;
  wire [0:0] wire_417;
  wire [0:0] wire_418;
  wire [63:0] wire_419;
  wire [0:0] wire_420;
  wire [31:0] wire_421;
  wire [7:0] wire_422;
  wire [0:0] wire_423;
  wire [63:0] wire_424;
  wire [0:0] wire_425;
  wire [0:0] wire_426;
  wire [63:0] wire_427;
  wire [0:0] wire_428;
  wire [31:0] wire_429;
  wire [31:0] wire_430;
  wire [7:0] wire_431;
  wire [31:0] wire_432;
  wire [7:0] wire_433;
  wire [0:0] wire_434;
  wire [7:0] wire_435;
  wire [31:0] wire_436;
  wire [7:0] wire_437;
  wire [0:0] wire_438;
  wire [7:0] wire_439;
  wire [0:0] wire_440;
  wire [0:0] wire_441;
  wire [0:0] wire_442;
  wire [7:0] wire_443;
  wire [31:0] wire_444;
  wire [7:0] wire_445;
  wire [0:0] wire_446;
  wire [0:0] wire_447;
  wire [31:0] wire_448;
  wire [0:0] wire_449;

endmodule
