module ALU (clk, rst, Register_1, Register_2, Instruction, Enable, PC, Error, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Register_1;
  input  wire [31:0] Register_2;
  input  wire [31:0] Instruction;
  input  wire [0:0] Enable;
  input  wire [31:0] PC;
  output  wire [0:0] Error;
  output  wire [31:0] Output;

  TC_Splitter32 # (.UUID(64'd856236723336969326 ^ UUID)) Splitter32_0 (.in(wire_25), .out0(wire_22), .out1(wire_81), .out2(), .out3(wire_73));
  TC_Splitter8 # (.UUID(64'd4590355626788055878 ^ UUID)) Splitter8_1 (.in(wire_22), .out0(), .out1(), .out2(wire_46), .out3(), .out4(), .out5(wire_6), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1157196835068389619 ^ UUID)) Splitter8_2 (.in(wire_73), .out0(), .out1(wire_2), .out2(wire_74), .out3(wire_51), .out4(wire_63), .out5(wire_17), .out6(wire_75), .out7());
  TC_Splitter8 # (.UUID(64'd2632572566828300203 ^ UUID)) Splitter8_3 (.in(wire_81), .out0(), .out1(), .out2(), .out3(), .out4(wire_84), .out5(wire_42), .out6(wire_24), .out7());
  TC_Switch # (.UUID(64'd2694834590265330456 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_4 (.en(wire_15), .in(wire_59), .out(wire_4_2));
  TC_Or # (.UUID(64'd1779458433257654647 ^ UUID), .BIT_WIDTH(64'd1)) Or_5 (.in0(wire_70), .in1(wire_56), .out(wire_82));
  TC_Or3 # (.UUID(64'd841580749221145212 ^ UUID), .BIT_WIDTH(64'd1)) Or3_6 (.in0(wire_74), .in1(wire_51), .in2(wire_63), .out(wire_110));
  TC_Or # (.UUID(64'd4480473029248294819 ^ UUID), .BIT_WIDTH(64'd1)) Or_7 (.in0(wire_110), .in1(wire_17), .out(wire_71));
  TC_Decoder3 # (.UUID(64'd1274385594707151563 ^ UUID)) Decoder3_8 (.dis(wire_91), .sel0(wire_84), .sel1(wire_42), .sel2(wire_24), .out0(wire_60), .out1(wire_32), .out2(wire_11), .out3(wire_67), .out4(wire_106), .out5(wire_0), .out6(wire_5), .out7(wire_86));
  TC_Mul # (.UUID(64'd426842451969131696 ^ UUID), .BIT_WIDTH(64'd32)) Mul32_9 (.in0(wire_29), .in1(wire_7), .out0(wire_72), .out1(wire_53));
  TC_Switch # (.UUID(64'd850462159983841261 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_10 (.en(wire_60), .in(wire_72), .out(wire_59_0));
  TC_Switch # (.UUID(64'd4359534044349454458 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_11 (.en(wire_32), .in(wire_53), .out(wire_59_1));
  TC_Switch # (.UUID(64'd1989058288848585541 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_12 (.en(wire_15), .in(wire_75), .out(wire_54));
  TC_Decoder3 # (.UUID(64'd1975167713134896394 ^ UUID)) Decoder3_13 (.dis(wire_87), .sel0(wire_84), .sel1(wire_42), .sel2(wire_24), .out0(wire_9), .out1(wire_47), .out2(wire_36), .out3(wire_39), .out4(wire_69), .out5(wire_38), .out6(wire_23), .out7(wire_76));
  TC_Not # (.UUID(64'd658721888043638227 ^ UUID), .BIT_WIDTH(64'd1)) Not_14 (.in(wire_31), .out(wire_87));
  TC_Not # (.UUID(64'd3401155971486664452 ^ UUID), .BIT_WIDTH(64'd1)) Not_15 (.in(wire_15), .out(wire_91));
  TC_Add # (.UUID(64'd4194481081827986572 ^ UUID), .BIT_WIDTH(64'd32)) Add32_16 (.in0(wire_29), .in1(wire_97), .ci(1'd0), .out(wire_37), .co());
  TC_Mux # (.UUID(64'd1954974504444484227 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_17 (.sel(wire_21), .in0(wire_12), .in1(wire_3), .out(wire_97));
  TC_Neg # (.UUID(64'd591805872178775221 ^ UUID), .BIT_WIDTH(64'd32)) Neg32_18 (.in(wire_12), .out(wire_3));
  TC_Switch # (.UUID(64'd462304321346859511 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_19 (.en(wire_9), .in(wire_37), .out(wire_1_5));
  TC_Switch # (.UUID(64'd4425345997042434399 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_20 (.en(wire_31), .in(wire_1), .out(wire_4_1));
  TC_Ashr # (.UUID(64'd3896657380015343184 ^ UUID), .BIT_WIDTH(64'd32)) Ashr32_21 (.in(wire_29), .shift(wire_12[7:0]), .out(wire_27));
  TC_Shl # (.UUID(64'd939190024179494840 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_22 (.in(wire_29), .shift(wire_12[7:0]), .out(wire_20));
  TC_Shr # (.UUID(64'd1111693115718089582 ^ UUID), .BIT_WIDTH(64'd32)) Shr32_23 (.in(wire_29), .shift(wire_12[7:0]), .out(wire_108));
  TC_Switch # (.UUID(64'd3021592203364150947 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_24 (.en(wire_47), .in(wire_20), .out(wire_1_3));
  TC_LessU # (.UUID(64'd2099414091277441902 ^ UUID), .BIT_WIDTH(64'd32)) LessU32_25 (.in0(wire_29), .in1(wire_12), .out(wire_57));
  TC_LessI # (.UUID(64'd359913812166468740 ^ UUID), .BIT_WIDTH(64'd32)) LessI32_26 (.in0(wire_29), .in1(wire_12), .out(wire_104));
  TC_Switch # (.UUID(64'd1156555378483579930 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_27 (.en(wire_36), .in({{31{1'b0}}, wire_104 }), .out(wire_1_0));
  TC_Switch # (.UUID(64'd2511188936079102141 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_28 (.en(wire_39), .in({{31{1'b0}}, wire_57 }), .out(wire_1_1));
  TC_Xor # (.UUID(64'd4070664494765303907 ^ UUID), .BIT_WIDTH(64'd32)) Xor32_29 (.in0(wire_29), .in1(wire_12), .out(wire_95));
  TC_Switch # (.UUID(64'd2710520328272254200 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_30 (.en(wire_69), .in(wire_95), .out(wire_1_2));
  TC_Switch # (.UUID(64'd2622542534940852509 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_31 (.en(wire_38), .in(wire_79), .out(wire_1_4));
  TC_Mux # (.UUID(64'd235825761551165049 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_32 (.sel(wire_21), .in0(wire_108), .in1(wire_27), .out(wire_79));
  TC_Or # (.UUID(64'd771507477978680572 ^ UUID), .BIT_WIDTH(64'd32)) Or32_33 (.in0(wire_29), .in1(wire_12), .out(wire_65));
  TC_And # (.UUID(64'd2644068751134878206 ^ UUID), .BIT_WIDTH(64'd32)) And32_34 (.in0(wire_29), .in1(wire_12), .out(wire_83));
  TC_Switch # (.UUID(64'd557390044361070583 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_35 (.en(wire_23), .in(wire_65), .out(wire_1_6));
  TC_Switch # (.UUID(64'd2699444628202921320 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_36 (.en(wire_76), .in(wire_83), .out(wire_1_7));
  TC_And # (.UUID(64'd695960843782682246 ^ UUID), .BIT_WIDTH(64'd1)) And_37 (.in0(wire_85), .in1(wire_71), .out(wire_56));
  TC_Or # (.UUID(64'd4262675205690804556 ^ UUID), .BIT_WIDTH(64'd1)) Or_38 (.in0(wire_19), .in1(wire_54), .out(wire_62));
  TC_Or # (.UUID(64'd1472109554877203089 ^ UUID), .BIT_WIDTH(64'd1)) Or_39 (.in0(wire_38), .in1(wire_47), .out(wire_109));
  TC_Mux # (.UUID(64'd3895625183492629013 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_40 (.sel(wire_6), .in0(wire_41), .in1(wire_7), .out(wire_12));
  TC_Switch # (.UUID(64'd4383360691348507301 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_15), .in(wire_6), .out(wire_112));
  TC_Or # (.UUID(64'd1190376895056596620 ^ UUID), .BIT_WIDTH(64'd1)) Or_42 (.in0(wire_62), .in1(wire_112), .out(wire_70));
  TC_And # (.UUID(64'd710606617466976572 ^ UUID), .BIT_WIDTH(64'd1)) And_43 (.in0(wire_48), .in1(wire_82), .out(wire_89));
  TC_Switch # (.UUID(64'd3384537657315157466 ^ UUID), .BIT_WIDTH(64'd32)) Output32z_44 (.en(wire_48), .in(wire_4), .out(Output));
  TC_Shr # (.UUID(64'd2917895975090633989 ^ UUID), .BIT_WIDTH(64'd32)) Shr32_45 (.in(wire_25), .shift(wire_64), .out());
  TC_Constant # (.UUID(64'd4133715739421574248 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h14)) Constant8_46 (.out(wire_64));
  TC_Shr # (.UUID(64'd1020156456611543410 ^ UUID), .BIT_WIDTH(64'd32)) Shr32_47 (.in(wire_25), .shift(wire_94), .out(wire_100));
  TC_Constant # (.UUID(64'd2865373584897540202 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h14)) Constant8_48 (.out(wire_94));
  TC_And # (.UUID(64'd485969331294057490 ^ UUID), .BIT_WIDTH(64'd8)) And8_49 (.in0(wire_100[7:0]), .in1(wire_92), .out(wire_50));
  TC_Constant # (.UUID(64'd2917838756477150323 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1F)) Constant8_50 (.out(wire_92));
  TC_Not # (.UUID(64'd547091731757834705 ^ UUID), .BIT_WIDTH(64'd1)) Not_51 (.in(wire_98), .out(wire_19));
  TC_Equal # (.UUID(64'd3672851681438596740 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_52 (.in0(wire_40), .in1(wire_80), .out(wire_98));
  TC_Constant # (.UUID(64'd25273916701498416 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h13)) Constant8_53 (.out(wire_40));
  TC_Maker8 # (.UUID(64'd3231735920723217485 ^ UUID)) Maker8_54 (.in0(wire_28), .in1(wire_102), .in2(1'd0), .in3(wire_105), .in4(wire_99), .in5(1'd0), .in6(wire_77), .in7(1'd0), .out(wire_80));
  TC_Splitter8 # (.UUID(64'd2624314861296391486 ^ UUID)) Splitter8_55 (.in(wire_22), .out0(wire_28), .out1(wire_102), .out2(), .out3(wire_105), .out4(wire_99), .out5(), .out6(wire_77), .out7());
  TC_And # (.UUID(64'd2124501545265996934 ^ UUID), .BIT_WIDTH(64'd1)) And_56 (.in0(wire_111), .in1(wire_49), .out(wire_31));
  TC_Not # (.UUID(64'd1806436245422777036 ^ UUID), .BIT_WIDTH(64'd1)) Not_57 (.in(wire_46), .out(wire_111));
  TC_And3 # (.UUID(64'd642894830652446579 ^ UUID), .BIT_WIDTH(64'd1)) And3_58 (.in0(wire_44), .in1(wire_6), .in2(wire_2), .out(wire_15));
  TC_Not # (.UUID(64'd2705641462022032447 ^ UUID), .BIT_WIDTH(64'd1)) Not_59 (.in(wire_46), .out(wire_44));
  TC_Switch # (.UUID(64'd1399457029941163327 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_60 (.en(wire_46), .in(wire_43), .out(wire_4_0));
  TC_Not # (.UUID(64'd248245287119840902 ^ UUID), .BIT_WIDTH(64'd1)) Not_61 (.in(wire_6), .out(wire_55));
  TC_Add # (.UUID(64'd4050497696309257697 ^ UUID), .BIT_WIDTH(64'd32)) Add32_62 (.in0(wire_33), .in1(wire_14), .ci(1'd0), .out(wire_16), .co());
  TC_Switch # (.UUID(64'd2971300873126547839 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_63 (.en(wire_55), .in(wire_16), .out(wire_43_0));
  TC_Constant # (.UUID(64'd312416627841680701 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFFFFF000)) Constant32_64 (.out(wire_8));
  TC_Switch # (.UUID(64'd3630921491077541815 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_65 (.en(wire_6), .in(wire_14), .out(wire_43_1));
  TC_And # (.UUID(64'd3522272529016663909 ^ UUID), .BIT_WIDTH(64'd32)) And32_66 (.in0(wire_25), .in1(wire_8), .out(wire_14));
  TC_Or # (.UUID(64'd2437551040465764240 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_113), .in1(wire_93), .out(wire_49));
  TC_Not # (.UUID(64'd4099482591278107694 ^ UUID), .BIT_WIDTH(64'd1)) Not_68 (.in(wire_6), .out(wire_113));
  TC_Not # (.UUID(64'd3939471549113845324 ^ UUID), .BIT_WIDTH(64'd1)) Not_69 (.in(wire_2), .out(wire_93));
  TC_And # (.UUID(64'd3857204907212449492 ^ UUID), .BIT_WIDTH(64'd1)) And_70 (.in0(wire_90), .in1(wire_6), .out(wire_85));
  TC_Not # (.UUID(64'd2156681183772808784 ^ UUID), .BIT_WIDTH(64'd1)) Not_71 (.in(wire_46), .out(wire_90));
  TC_Splitter8 # (.UUID(64'd4290930814921900217 ^ UUID)) Splitter8_72 (.in(wire_45), .out0(wire_35), .out1(wire_68), .out2(wire_107), .out3(wire_66), .out4(wire_34), .out5(wire_88), .out6(wire_78), .out7(wire_13));
  TC_Maker8 # (.UUID(64'd4186148599523492260 ^ UUID)) Maker8_73 (.in0(wire_34), .in1(wire_88), .in2(wire_78), .in3(wire_13), .in4(wire_13), .in5(wire_13), .in6(wire_13), .in7(wire_13), .out(wire_18));
  TC_Maker8 # (.UUID(64'd1075353434363615074 ^ UUID)) Maker8_74 (.in0(wire_13), .in1(wire_13), .in2(wire_13), .in3(wire_13), .in4(wire_13), .in5(wire_13), .in6(wire_13), .in7(wire_13), .out(wire_10));
  TC_Maker8 # (.UUID(64'd1323227554668416689 ^ UUID)) Maker8_75 (.in0(wire_13), .in1(wire_13), .in2(wire_13), .in3(wire_13), .in4(wire_13), .in5(wire_13), .in6(wire_13), .in7(wire_13), .out(wire_58));
  TC_Maker8 # (.UUID(64'd1235368889047368006 ^ UUID)) Maker8_76 (.in0(wire_103), .in1(wire_61), .in2(wire_101), .in3(wire_26), .in4(wire_35), .in5(wire_68), .in6(wire_107), .in7(wire_66), .out(wire_96));
  TC_Splitter8 # (.UUID(64'd3679310397701514836 ^ UUID)) Splitter8_77 (.in(wire_52), .out0(), .out1(), .out2(), .out3(), .out4(wire_103), .out5(wire_61), .out6(wire_101), .out7(wire_26));
  TC_Splitter32 # (.UUID(64'd740850826075132075 ^ UUID)) Splitter32_78 (.in(wire_25), .out0(), .out1(), .out2(wire_52), .out3(wire_45));
  TC_Maker32 # (.UUID(64'd408416054360199427 ^ UUID)) Maker32_79 (.in0(wire_96), .in1(wire_18), .in2(wire_10), .in3(wire_58), .out(wire_30));
  TC_Mux # (.UUID(64'd3673667422785486178 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_80 (.sel(wire_109), .in0(wire_30), .in1({{24{1'b0}}, wire_50 }), .out(wire_41));
  TC_And # (.UUID(64'd53600999146838859 ^ UUID), .BIT_WIDTH(64'd1)) And_81 (.in0(wire_75), .in1(wire_6), .out(wire_21));

  wire [0:0] wire_0;
  wire [31:0] wire_1;
  wire [31:0] wire_1_0;
  wire [31:0] wire_1_1;
  wire [31:0] wire_1_2;
  wire [31:0] wire_1_3;
  wire [31:0] wire_1_4;
  wire [31:0] wire_1_5;
  wire [31:0] wire_1_6;
  wire [31:0] wire_1_7;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7;
  wire [0:0] wire_2;
  wire [31:0] wire_3;
  wire [31:0] wire_4;
  wire [31:0] wire_4_0;
  wire [31:0] wire_4_1;
  wire [31:0] wire_4_2;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [31:0] wire_7;
  assign wire_7 = Register_2;
  wire [31:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [31:0] wire_12;
  wire [0:0] wire_13;
  wire [31:0] wire_14;
  wire [0:0] wire_15;
  wire [31:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [31:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [31:0] wire_25;
  assign wire_25 = Instruction;
  wire [0:0] wire_26;
  wire [31:0] wire_27;
  wire [0:0] wire_28;
  wire [31:0] wire_29;
  assign wire_29 = Register_1;
  wire [31:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [31:0] wire_33;
  assign wire_33 = PC;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [31:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [31:0] wire_41;
  wire [0:0] wire_42;
  wire [31:0] wire_43;
  wire [31:0] wire_43_0;
  wire [31:0] wire_43_1;
  assign wire_43 = wire_43_0|wire_43_1;
  wire [0:0] wire_44;
  wire [7:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  assign wire_48 = Enable;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [31:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [31:0] wire_59;
  wire [31:0] wire_59_0;
  wire [31:0] wire_59_1;
  assign wire_59 = wire_59_0|wire_59_1;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [7:0] wire_64;
  wire [31:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [31:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [31:0] wire_79;
  wire [7:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [31:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  assign Error = wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [7:0] wire_92;
  wire [0:0] wire_93;
  wire [7:0] wire_94;
  wire [31:0] wire_95;
  wire [7:0] wire_96;
  wire [31:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [31:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [31:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;

endmodule
