module LEG_ALU (clk, rst, \�_____ , \�______1 , \�______2 , Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] \�_____ ;
  input  wire [7:0] \�______1 ;
  input  wire [7:0] \�______2 ;
  output  wire [7:0] Output;

  TC_Splitter8 # (.UUID(64'd4503754288184316976 ^ UUID)) Splitter8_0 (.in(wire_15), .out0(wire_30), .out1(wire_8), .out2(wire_28), .out3(wire_5), .out4(), .out5(), .out6(), .out7());
  TC_Or # (.UUID(64'd2102355290693069281 ^ UUID), .BIT_WIDTH(64'd8)) Or8_1 (.in0(wire_1), .in1(wire_2), .out(wire_26));
  TC_Switch # (.UUID(64'd3955843348845505503 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_2 (.en(wire_6), .in(wire_26), .out(wire_3_0));
  TC_Or # (.UUID(64'd1138358230590770772 ^ UUID), .BIT_WIDTH(64'd8)) Or8_3 (.in0(wire_12), .in1(wire_17), .out(wire_18));
  TC_Not # (.UUID(64'd2874953002594435817 ^ UUID), .BIT_WIDTH(64'd8)) Not8_4 (.in(wire_1), .out(wire_12));
  TC_Not # (.UUID(64'd3261420662032331478 ^ UUID), .BIT_WIDTH(64'd8)) Not8_5 (.in(wire_2), .out(wire_17));
  TC_Switch # (.UUID(64'd1559193756622028187 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_24), .in(wire_18), .out(wire_3_3));
  TC_Switch # (.UUID(64'd562902586904156559 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_13), .in(wire_9), .out(wire_3_2));
  TC_Or # (.UUID(64'd1762851381222581582 ^ UUID), .BIT_WIDTH(64'd8)) Or8_8 (.in0(wire_1), .in1(wire_2), .out(wire_19));
  TC_Not # (.UUID(64'd3866306404953024228 ^ UUID), .BIT_WIDTH(64'd8)) Not8_9 (.in(wire_19), .out(wire_9));
  TC_Not # (.UUID(64'd4374362103234097039 ^ UUID), .BIT_WIDTH(64'd8)) Not8_10 (.in(wire_1), .out(wire_16));
  TC_Not # (.UUID(64'd1299975577945567859 ^ UUID), .BIT_WIDTH(64'd8)) Not8_11 (.in(wire_2), .out(wire_0));
  TC_Or # (.UUID(64'd3778950935273956021 ^ UUID), .BIT_WIDTH(64'd8)) Or8_12 (.in0(wire_16), .in1(wire_0), .out(wire_23));
  TC_Not # (.UUID(64'd1920809211267629108 ^ UUID), .BIT_WIDTH(64'd8)) Not8_13 (.in(wire_23), .out(wire_27));
  TC_Switch # (.UUID(64'd3823930859173339200 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_7), .in(wire_27), .out(wire_3_1));
  TC_Switch # (.UUID(64'd3202039647240155243 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_29), .in(wire_21), .out(wire_3_4));
  TC_Add # (.UUID(64'd2569020168253982736 ^ UUID), .BIT_WIDTH(64'd8)) Add8_16 (.in0(wire_1), .in1(wire_2), .ci(1'd0), .out(wire_21), .co());
  TC_Switch # (.UUID(64'd2734422171326569155 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_4), .in(wire_25), .out(wire_3_7));
  TC_Add # (.UUID(64'd4595643146173721565 ^ UUID), .BIT_WIDTH(64'd8)) Add8_18 (.in0(wire_1), .in1(wire_11), .ci(1'd0), .out(wire_25), .co());
  TC_Neg # (.UUID(64'd4435798358922345065 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_19 (.in(wire_2), .out(wire_11));
  _4bit_Decoder # (.UUID(64'd1725263961771509634 ^ UUID)) _4bit_Decoder_20 (.clk(clk), .rst(rst), .\1_1 (wire_30), .\2_1 (wire_8), .\4_1 (wire_28), .\8_1 (wire_5), .\7 (), .\11 (), .\3 (wire_6), .\15 (wire_24), .\6 (), .\8_2 (), .\5 (wire_20), .\9 (), .\10 (), .\4_2 (wire_22), .\12 (), .\13 (), .\14 (wire_13), .\2_2 (wire_7), .\1_2 (wire_4), .\0 (wire_29));
  TC_Switch # (.UUID(64'd1852877134885786992 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_22), .in(wire_10), .out(wire_3_5));
  TC_Not # (.UUID(64'd2650145618189716223 ^ UUID), .BIT_WIDTH(64'd8)) Not8_22 (.in(wire_1), .out(wire_10));
  TC_Xor # (.UUID(64'd457105424950704873 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_23 (.in0(wire_1), .in1(wire_2), .out(wire_14));
  TC_Switch # (.UUID(64'd2882176525213117412 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_20), .in(wire_14), .out(wire_3_6));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  assign wire_1 = \�______1 ;
  wire [7:0] wire_2;
  assign wire_2 = \�______2 ;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7;
  assign Output = wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [7:0] wire_15;
  assign wire_15 = \�_____ ;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;

endmodule
