module Controlz_Block (clk, rst, Instruction, Register_1, Register_2, Enabled, PC, Register_Out, Write_Register, PC_Out, Should_Jump);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Instruction;
  input  wire [31:0] Register_1;
  input  wire [31:0] Register_2;
  input  wire [0:0] Enabled;
  input  wire [31:0] PC;
  output  wire [31:0] Register_Out;
  output  wire [0:0] Write_Register;
  output  wire [31:0] PC_Out;
  output  wire [0:0] Should_Jump;

  TC_Splitter8 # (.UUID(64'd902104352047372224 ^ UUID)) Splitter8_0 (.in(wire_43), .out0(), .out1(), .out2(wire_40), .out3(wire_37), .out4(), .out5(), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd1707422630313500119 ^ UUID)) Splitter32_1 (.in(wire_11), .out0(wire_43), .out1(wire_63), .out2(), .out3());
  TC_Switch # (.UUID(64'd1996006586573775508 ^ UUID), .BIT_WIDTH(64'd32)) Output32z_2 (.en(wire_27), .in(wire_2), .out(PC_Out));
  TC_Splitter8 # (.UUID(64'd3577095691572030781 ^ UUID)) Splitter8_3 (.in(wire_63), .out0(), .out1(), .out2(), .out3(), .out4(wire_13), .out5(wire_65), .out6(wire_14), .out7());
  TC_And # (.UUID(64'd3038231527070571591 ^ UUID), .BIT_WIDTH(64'd1)) And_4 (.in0(wire_27), .in1(wire_87), .out(wire_92));
  TC_Not # (.UUID(64'd1823206584575818658 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_40), .out(wire_4));
  TC_Decoder3 # (.UUID(64'd687181082384468536 ^ UUID)) Decoder3_6 (.dis(wire_24), .sel0(wire_13), .sel1(wire_65), .sel2(wire_14), .out0(wire_61), .out1(wire_76), .out2(wire_20), .out3(wire_62), .out4(wire_47), .out5(wire_9), .out6(wire_12), .out7(wire_28));
  TC_Equal # (.UUID(64'd2633171923279527042 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_7 (.in0(wire_34), .in1(wire_6), .out(wire_48));
  TC_Add # (.UUID(64'd4517514505079768302 ^ UUID), .BIT_WIDTH(64'd32)) Add32_8 (.in0(wire_55), .in1(wire_57), .ci(1'd0), .out(wire_72), .co());
  TC_Switch # (.UUID(64'd1337027801841510438 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_9 (.en(wire_4), .in(wire_72), .out(wire_2_1));
  TC_Switch # (.UUID(64'd79888115093657123 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_10 (.en(wire_61), .in(wire_48), .out(wire_15_5));
  TC_Switch # (.UUID(64'd3274754959937476190 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_76), .in(wire_44), .out(wire_15_4));
  TC_Not # (.UUID(64'd4395154833012517612 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_48), .out(wire_44));
  TC_Switch # (.UUID(64'd4399928849220487887 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_13 (.en(wire_4), .in(wire_15), .out(wire_22));
  TC_LessI # (.UUID(64'd2922862214185537558 ^ UUID), .BIT_WIDTH(64'd32)) LessI32_14 (.in0(wire_34), .in1(wire_6), .out(wire_95));
  TC_LessU # (.UUID(64'd1879850586635247184 ^ UUID), .BIT_WIDTH(64'd32)) LessU32_15 (.in0(wire_34), .in1(wire_6), .out(wire_25));
  TC_Switch # (.UUID(64'd4203613056368251062 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_16 (.en(wire_47), .in(wire_95), .out(wire_15_3));
  TC_Switch # (.UUID(64'd4548650618125891994 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_12), .in(wire_25), .out(wire_15_0));
  TC_Switch # (.UUID(64'd3895235215987418618 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_9), .in(wire_77), .out(wire_15_2));
  TC_Switch # (.UUID(64'd3867017945406718342 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_19 (.en(wire_28), .in(wire_78), .out(wire_15_1));
  TC_Not # (.UUID(64'd1084624806982300785 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_95), .out(wire_77));
  TC_Not # (.UUID(64'd2960215855915062300 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_25), .out(wire_78));
  TC_Not # (.UUID(64'd2873907438454793039 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_4), .out(wire_24));
  TC_And # (.UUID(64'd1529293667396716322 ^ UUID), .BIT_WIDTH(64'd1)) And_23 (.in0(wire_27), .in1(wire_40), .out(wire_108));
  TC_Splitter8 # (.UUID(64'd4515631532377864634 ^ UUID)) Splitter8_24 (.in(wire_30), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_103));
  TC_Splitter8 # (.UUID(64'd4078659507003827988 ^ UUID)) Splitter8_25 (.in(wire_84), .out0(wire_53), .out1(wire_91), .out2(wire_93), .out3(wire_60), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2134980236709436119 ^ UUID)) Splitter8_26 (.in(wire_21), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2952686544166958164 ^ UUID)) Splitter8_27 (.in(wire_5), .out0(), .out1(wire_36), .out2(wire_46), .out3(wire_54), .out4(wire_89), .out5(wire_42), .out6(wire_51), .out7(wire_0));
  TC_Maker8 # (.UUID(64'd2008199746892869203 ^ UUID)) Maker8_28 (.in0(wire_0), .in1(wire_0), .in2(wire_0), .in3(wire_0), .in4(wire_0), .in5(wire_0), .in6(wire_0), .in7(wire_0), .out(wire_99));
  TC_Maker8 # (.UUID(64'd4590122625182198597 ^ UUID)) Maker8_29 (.in0(wire_0), .in1(wire_0), .in2(wire_0), .in3(wire_0), .in4(wire_0), .in5(wire_0), .in6(wire_0), .in7(wire_0), .out(wire_80));
  TC_Maker8 # (.UUID(64'd610578434292512677 ^ UUID)) Maker8_30 (.in0(wire_89), .in1(wire_42), .in2(wire_51), .in3(wire_103), .in4(wire_0), .in5(wire_0), .in6(wire_0), .in7(wire_0), .out(wire_69));
  TC_Maker8 # (.UUID(64'd2852305094401698312 ^ UUID)) Maker8_31 (.in0(1'd0), .in1(wire_53), .in2(wire_91), .in3(wire_93), .in4(wire_60), .in5(wire_36), .in6(wire_46), .in7(wire_54), .out(wire_73));
  TC_Maker32 # (.UUID(64'd241392417761818401 ^ UUID)) Maker32_32 (.in0(wire_73), .in1(wire_69), .in2(wire_80), .in3(wire_99), .out(wire_55));
  TC_Splitter32 # (.UUID(64'd647400026824596760 ^ UUID)) Splitter32_33 (.in(wire_11), .out0(wire_30), .out1(wire_84), .out2(wire_21), .out3(wire_5));
  TC_And # (.UUID(64'd981401743066463860 ^ UUID), .BIT_WIDTH(64'd1)) And_34 (.in0(wire_37), .in1(wire_40), .out(wire_85));
  TC_Splitter32 # (.UUID(64'd2678735073178107162 ^ UUID)) Splitter32_35 (.in(wire_11), .out0(), .out1(wire_31), .out2(wire_29), .out3(wire_75));
  TC_Splitter8 # (.UUID(64'd2335251480870319275 ^ UUID)) Splitter8_36 (.in(wire_31), .out0(), .out1(), .out2(), .out3(), .out4(wire_58), .out5(wire_105), .out6(wire_71), .out7(wire_86));
  TC_Splitter8 # (.UUID(64'd1559009683295488391 ^ UUID)) Splitter8_37 (.in(wire_29), .out0(wire_106), .out1(wire_33), .out2(wire_67), .out3(wire_19), .out4(wire_16), .out5(wire_94), .out6(wire_101), .out7(wire_41));
  TC_Splitter8 # (.UUID(64'd4227780176090406672 ^ UUID)) Splitter8_38 (.in(wire_75), .out0(wire_109), .out1(wire_45), .out2(wire_100), .out3(wire_64), .out4(wire_107), .out5(wire_70), .out6(wire_49), .out7(wire_32));
  TC_Maker8 # (.UUID(64'd2878091998981806722 ^ UUID)) Maker8_39 (.in0(1'd0), .in1(wire_94), .in2(wire_101), .in3(wire_41), .in4(wire_109), .in5(wire_45), .in6(wire_100), .in7(wire_64), .out(wire_10));
  TC_Maker32 # (.UUID(64'd2407390854939498277 ^ UUID)) Maker32_40 (.in0(wire_10), .in1(wire_97), .in2(wire_52), .in3(wire_8), .out(wire_79));
  TC_Maker8 # (.UUID(64'd301639447571383139 ^ UUID)) Maker8_41 (.in0(wire_107), .in1(wire_70), .in2(wire_49), .in3(wire_16), .in4(wire_58), .in5(wire_105), .in6(wire_71), .in7(wire_86), .out(wire_97));
  TC_Maker8 # (.UUID(64'd3387325518231762438 ^ UUID)) Maker8_42 (.in0(wire_106), .in1(wire_33), .in2(wire_67), .in3(wire_19), .in4(wire_32), .in5(wire_32), .in6(wire_32), .in7(wire_32), .out(wire_52));
  TC_Maker8 # (.UUID(64'd88120391011758893 ^ UUID)) Maker8_43 (.in0(wire_32), .in1(wire_32), .in2(wire_32), .in3(wire_32), .in4(wire_32), .in5(wire_32), .in6(wire_32), .in7(wire_32), .out(wire_8));
  TC_Switch # (.UUID(64'd3456175386122381956 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_44 (.en(wire_85), .in(wire_23), .out(wire_2_0));
  TC_And # (.UUID(64'd4143119125227311513 ^ UUID), .BIT_WIDTH(64'd1)) And_45 (.in0(wire_1), .in1(wire_40), .out(wire_35));
  TC_Not # (.UUID(64'd2111987689116572799 ^ UUID), .BIT_WIDTH(64'd1)) Not_46 (.in(wire_37), .out(wire_1));
  TC_Switch # (.UUID(64'd270105768238044738 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_47 (.en(wire_35), .in(wire_50), .out(wire_2_2));
  TC_Add # (.UUID(64'd4320218808739467258 ^ UUID), .BIT_WIDTH(64'd32)) Add32_48 (.in0(wire_34), .in1(wire_59), .ci(1'd0), .out(wire_68), .co());
  TC_Splitter32 # (.UUID(64'd821229586171559223 ^ UUID)) Splitter32_49 (.in(wire_11), .out0(), .out1(), .out2(wire_38), .out3(wire_3));
  TC_Splitter8 # (.UUID(64'd2728032006665629024 ^ UUID)) Splitter8_50 (.in(wire_38), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(wire_26), .out6(wire_110), .out7(wire_66));
  TC_Splitter8 # (.UUID(64'd3065001218220038661 ^ UUID)) Splitter8_51 (.in(wire_3), .out0(wire_88), .out1(wire_82), .out2(wire_90), .out3(wire_104), .out4(wire_102), .out5(wire_17), .out6(wire_98), .out7(wire_18));
  TC_Maker8 # (.UUID(64'd2989533700026571770 ^ UUID)) Maker8_52 (.in0(1'd0), .in1(wire_26), .in2(wire_110), .in3(wire_66), .in4(wire_88), .in5(wire_82), .in6(wire_90), .in7(wire_104), .out(wire_39));
  TC_Maker8 # (.UUID(64'd2542130407660439527 ^ UUID)) Maker8_53 (.in0(wire_102), .in1(wire_17), .in2(wire_98), .in3(wire_18), .in4(wire_18), .in5(wire_18), .in6(wire_18), .in7(wire_18), .out(wire_7));
  TC_Maker32 # (.UUID(64'd1044328868542777178 ^ UUID)) Maker32_54 (.in0(wire_39), .in1(wire_7), .in2(wire_56), .in3(wire_81), .out(wire_59));
  TC_And # (.UUID(64'd2761644439738323318 ^ UUID), .BIT_WIDTH(64'd32)) And32_55 (.in0(wire_68), .in1(wire_74), .out(wire_50));
  TC_Constant # (.UUID(64'd2839113499863336469 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFFFFFFFE)) Constant32_56 (.out(wire_74));
  TC_Or # (.UUID(64'd2052510646991599899 ^ UUID), .BIT_WIDTH(64'd1)) Or_57 (.in0(wire_22), .in1(wire_40), .out(wire_87));
  TC_Switch # (.UUID(64'd1041243192545914942 ^ UUID), .BIT_WIDTH(64'd32)) Output32z_58 (.en(wire_27), .in(wire_83), .out(Register_Out));
  TC_Add # (.UUID(64'd4227437673484616104 ^ UUID), .BIT_WIDTH(64'd32)) Add32_59 (.in0(wire_57), .in1({{24{1'b0}}, wire_96 }), .ci(1'd0), .out(wire_83), .co());
  TC_Constant # (.UUID(64'd1872495430187045921 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_60 (.out(wire_96));
  TC_Add # (.UUID(64'd4034940777489028077 ^ UUID), .BIT_WIDTH(64'd32)) Add32_61 (.in0(wire_57), .in1(wire_79), .ci(1'd0), .out(wire_23), .co());
  TC_Maker8 # (.UUID(64'd4042000985687822218 ^ UUID)) Maker8_62 (.in0(wire_18), .in1(wire_18), .in2(wire_18), .in3(wire_18), .in4(wire_18), .in5(wire_18), .in6(wire_18), .in7(wire_18), .out(wire_56));
  TC_Maker8 # (.UUID(64'd3617674189833292210 ^ UUID)) Maker8_63 (.in0(wire_18), .in1(wire_18), .in2(wire_18), .in3(wire_18), .in4(wire_18), .in5(wire_18), .in6(wire_18), .in7(wire_18), .out(wire_81));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [31:0] wire_2;
  wire [31:0] wire_2_0;
  wire [31:0] wire_2_1;
  wire [31:0] wire_2_2;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [31:0] wire_6;
  assign wire_6 = Register_2;
  wire [7:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [31:0] wire_11;
  assign wire_11 = Instruction;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_15_0;
  wire [0:0] wire_15_1;
  wire [0:0] wire_15_2;
  wire [0:0] wire_15_3;
  wire [0:0] wire_15_4;
  wire [0:0] wire_15_5;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3|wire_15_4|wire_15_5;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [31:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  assign wire_27 = Enabled;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [31:0] wire_34;
  assign wire_34 = Register_1;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [31:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [31:0] wire_55;
  wire [7:0] wire_56;
  wire [31:0] wire_57;
  assign wire_57 = PC;
  wire [0:0] wire_58;
  wire [31:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [31:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [31:0] wire_72;
  wire [7:0] wire_73;
  wire [31:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [31:0] wire_79;
  wire [7:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [31:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  assign Should_Jump = wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [7:0] wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [7:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  assign Write_Register = wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;

endmodule
