module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_3), .en(wire_9), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_93), .in(arch_input_value), .out(wire_12));
  TC_Counter # (.UUID(64'd1175999672554394000 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_2 (.clk(clk), .rst(rst), .save(wire_64), .in(wire_3), .out(wire_35));
  TC_Splitter8 # (.UUID(64'd3496280010280654809 ^ UUID)) Splitter8_3 (.in(wire_15), .out0(wire_95), .out1(wire_60), .out2(wire_105), .out3(wire_40), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1350359362790102949 ^ UUID)) Splitter8_4 (.in(wire_81), .out0(wire_85), .out1(wire_42), .out2(wire_6), .out3(wire_104), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3688384451292696869 ^ UUID)) Splitter8_5 (.in(wire_53), .out0(wire_102), .out1(wire_86), .out2(wire_62), .out3(wire_103), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3357720912797461292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_77), .in(wire_35), .out());
  TC_Maker8 # (.UUID(64'd2922775923237819214 ^ UUID)) Maker8_7 (.in0(wire_88), .in1(wire_61), .in2(wire_34), .in3(wire_97), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_58));
  TC_Splitter8 # (.UUID(64'd4136660363423911410 ^ UUID)) Splitter8_8 (.in(wire_8[7:0]), .out0(wire_88), .out1(wire_61), .out2(wire_34), .out3(wire_97), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd4550958897663313502 ^ UUID)) Splitter8_9 (.in(wire_8[7:0]), .out0(wire_67), .out1(wire_26), .out2(wire_24), .out3(wire_78), .out4(wire_107), .out5(wire_66), .out6(wire_115), .out7(wire_89));
  TC_Maker8 # (.UUID(64'd3153840370766490713 ^ UUID)) Maker8_10 (.in0(wire_67), .in1(wire_26), .in2(wire_24), .in3(wire_78), .in4(wire_107), .in5(wire_66), .in6(wire_115), .in7(wire_89), .out(wire_4));
  TC_Constant # (.UUID(64'd4029987529778329422 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out(wire_96));
  TC_Constant # (.UUID(64'd47372170638122597 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out(wire_33));
  TC_Constant # (.UUID(64'd3010400910295959985 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_80));
  TC_Constant # (.UUID(64'd1353887318054096472 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_109));
  TC_Constant # (.UUID(64'd4461919415197064488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out(wire_94));
  TC_Constant # (.UUID(64'd2551986311311524963 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_108));
  TC_Switch # (.UUID(64'd201407107924193690 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_118), .in(wire_44), .out(wire_0_1));
  TC_Switch # (.UUID(64'd3784926049681585699 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_75), .in(wire_44), .out(wire_10_6));
  TC_Switch # (.UUID(64'd3418942253385023549 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_83), .in(wire_11), .out(wire_0_6));
  TC_Switch # (.UUID(64'd3104771108315787100 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_65), .in(wire_11), .out(wire_10_4));
  TC_Switch # (.UUID(64'd494263610589549334 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_51), .in(wire_28), .out(wire_0_0));
  TC_Switch # (.UUID(64'd4455028313033582898 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_59), .in(wire_28), .out(wire_10_3));
  TC_Switch # (.UUID(64'd977062972681925203 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_90), .in(wire_41), .out(wire_0_4));
  TC_Switch # (.UUID(64'd2935373336597064260 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_32), .in(wire_41), .out(wire_10_1));
  TC_Switch # (.UUID(64'd2595310988575568445 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_52), .in(wire_46), .out(wire_0_3));
  TC_Switch # (.UUID(64'd3649926646471230167 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_87), .in(wire_46), .out(wire_10_5));
  TC_Switch # (.UUID(64'd115863760055946247 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_25), .in(wire_39), .out(wire_0_2));
  TC_Switch # (.UUID(64'd459043271910661458 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_20), .in(wire_39), .out(wire_10_2));
  TC_Switch # (.UUID(64'd4275937720180353902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_114), .in(wire_35), .out());
  TC_Switch # (.UUID(64'd2718446434835356700 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_54), .in(wire_12), .out(wire_0_5));
  TC_Switch # (.UUID(64'd1811299859375739998 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_17), .in(wire_12), .out(wire_10_0));
  TC_Or # (.UUID(64'd117421755651659184 ^ UUID), .BIT_WIDTH(64'd1)) Or_32 (.in0(wire_54), .in1(wire_17), .out(wire_93));
  TC_Switch # (.UUID(64'd262409980643160938 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_49), .in(wire_45[7:0]), .out(wire_10_10));
  TC_Switch # (.UUID(64'd2764614579549035605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_56), .in(wire_73[7:0]), .out(wire_0_8));
  TC_Switch # (.UUID(64'd2974460371787013801 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_113), .in(wire_111), .out(wire_3_0));
  TC_Mux # (.UUID(64'd1769789085559769130 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_36 (.sel(wire_49), .in0(wire_45[7:0]), .in1(wire_21), .out(wire_81));
  TC_Mux # (.UUID(64'd1404337327044278632 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_37 (.sel(wire_56), .in0(wire_73[7:0]), .in1(wire_98), .out(wire_15));
  TC_Constant # (.UUID(64'd4387708643330744374 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_38 (.out(wire_98));
  TC_Constant # (.UUID(64'd2430039925245603401 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_39 (.out(wire_21));
  TC_Switch # (.UUID(64'd3877536405880520929 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_92), .in(wire_69), .out(wire_36));
  TC_Constant # (.UUID(64'd2430392602802046886 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_41 (.out(wire_57));
  TC_Mux # (.UUID(64'd1559488034901936773 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_42 (.sel(wire_36), .in0(wire_91), .in1(wire_57), .out(wire_53));
  TC_Switch # (.UUID(64'd3981948550050450551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_36), .in(wire_19[7:0]), .out(wire_3_1));
  TC_Ram # (.UUID(64'd1683242105781375453 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_44 (.clk(clk), .rst(rst), .load(wire_68), .save(wire_18), .address({{24{1'b0}}, wire_82 }), .in0({{56{1'b0}}, wire_3 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_16), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd1949247607308932292 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_45 (.out(wire_84));
  TC_Or # (.UUID(64'd2571069615494455195 ^ UUID), .BIT_WIDTH(64'd1)) Or_46 (.in0(wire_47), .in1(wire_23), .out(wire_68));
  TC_Switch # (.UUID(64'd3896516251333244950 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_48), .in(wire_14), .out(wire_0_7));
  TC_Switch # (.UUID(64'd4219278115069450234 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_5), .in(wire_14), .out(wire_10_7));
  TC_Switch # (.UUID(64'd875265095609107539 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_47), .in(wire_16[7:0]), .out(wire_0_10));
  TC_Switch # (.UUID(64'd1025433274855748469 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_23), .in(wire_16[7:0]), .out(wire_10_8));
  TC_Program # (.UUID(64'd4489305393227859486 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_3E4D37784397861E.w8.bin"), .ARG_SIG("Program_3E4D37784397861E=%s")) Program_51 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_35 }), .out0(wire_8), .out1(wire_73), .out2(wire_45), .out3(wire_19));
  TC_Switch # (.UUID(64'd3036050060892365836 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_74), .in(wire_38), .out(wire_0_9));
  TC_Switch # (.UUID(64'd3830579770898048556 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_1), .in(wire_38), .out(wire_10_9));
  TC_Or # (.UUID(64'd1511395350716789461 ^ UUID), .BIT_WIDTH(64'd1)) Or_54 (.in0(wire_74), .in1(wire_1), .out(wire_31));
  _4bit_Decoder # (.UUID(64'd188593635878702660 ^ UUID)) _4bit_Decoder_55 (.clk(clk), .rst(rst), .\1_1 (wire_95), .\2_1 (wire_60), .\4_1 (wire_105), .\8_1 (wire_40), .\7 (wire_54), .\11 (), .\3 (wire_90), .\15 (), .\6 (wire_77), .\8_2 (wire_48), .\5 (wire_25), .\9 (wire_47), .\10 (wire_74), .\4_2 (wire_52), .\12 (), .\13 (), .\14 (), .\2_2 (wire_51), .\1_2 (wire_83), .\0 (wire_118));
  _4bit_Decoder # (.UUID(64'd3657203059375966986 ^ UUID)) _4bit_Decoder_56 (.clk(clk), .rst(rst), .\1_1 (wire_85), .\2_1 (wire_42), .\4_1 (wire_6), .\8_1 (wire_104), .\7 (wire_17), .\11 (), .\3 (wire_32), .\15 (), .\6 (wire_114), .\8_2 (wire_5), .\5 (wire_20), .\9 (wire_23), .\10 (wire_1), .\4_2 (wire_87), .\12 (), .\13 (), .\14 (), .\2_2 (wire_59), .\1_2 (wire_65), .\0 (wire_75));
  _4bit_Decoder # (.UUID(64'd4526675728054865805 ^ UUID)) _4bit_Decoder_57 (.clk(clk), .rst(rst), .\1_1 (wire_102), .\2_1 (wire_86), .\4_1 (wire_62), .\8_1 (wire_103), .\7 (wire_9), .\11 (), .\3 (wire_50), .\15 (), .\6 (wire_64), .\8_2 (wire_27), .\5 (wire_79), .\9 (wire_18), .\10 (wire_30), .\4_2 (wire_117), .\12 (), .\13 (), .\14 (), .\2_2 (wire_71), .\1_2 (wire_70), .\0 (wire_116));
  RegisterPlus # (.UUID(64'd1898575026262245003 ^ UUID)) RegisterPlus_58 (.clk(clk), .rst(rst), .\�_____ (wire_96), .\�___________ (wire_3), .\�_____ (wire_116), .\�___________ (), .Output(wire_44));
  RegisterPlus # (.UUID(64'd201486149512558618 ^ UUID)) RegisterPlus_59 (.clk(clk), .rst(rst), .\�_____ (wire_33), .\�___________ (wire_3), .\�_____ (wire_70), .\�___________ (), .Output(wire_11));
  RegisterPlus # (.UUID(64'd4130910523704063521 ^ UUID)) RegisterPlus_60 (.clk(clk), .rst(rst), .\�_____ (wire_80), .\�___________ (wire_3), .\�_____ (wire_71), .\�___________ (), .Output(wire_28));
  RegisterPlus # (.UUID(64'd579904311903668382 ^ UUID)) RegisterPlus_61 (.clk(clk), .rst(rst), .\�_____ (wire_109), .\�___________ (wire_3), .\�_____ (wire_50), .\�___________ (), .Output(wire_41));
  RegisterPlus # (.UUID(64'd2026589517635316452 ^ UUID)) RegisterPlus_62 (.clk(clk), .rst(rst), .\�_____ (wire_94), .\�___________ (wire_3), .\�_____ (wire_117), .\�___________ (), .Output(wire_46));
  RegisterPlus # (.UUID(64'd1622410096212380183 ^ UUID)) RegisterPlus_63 (.clk(clk), .rst(rst), .\�_____ (wire_108), .\�___________ (wire_3), .\�_____ (wire_79), .\�___________ (), .Output(wire_39));
  LEG_COND # (.UUID(64'd999600516743479399 ^ UUID)) LEG_COND_64 (.clk(clk), .rst(rst), .ARG1(wire_0), .ARG2(wire_10), .\�_____ (wire_8[7:0]), .Output(wire_69));
  RegisterPlus # (.UUID(64'd471658098348471390 ^ UUID)) RegisterPlus_65 (.clk(clk), .rst(rst), .\�_____ (wire_84), .\�___________ (wire_3), .\�_____ (wire_27), .\�___________ (wire_82), .Output(wire_14));
  LEG_DEC # (.UUID(64'd2015393024950033718 ^ UUID)) LEG_DEC_66 (.clk(clk), .rst(rst), .OPCODE(wire_4), .IMMEDIATE1(wire_56), .IMMEDIATE2(wire_49), .CALCULATION(wire_113), .JUMP(wire_92));
  ZXE6ZXA0ZX88 # (.UUID(64'd1806005441980126369 ^ UUID)) ZXE6ZXA0ZX88_67 (.clk(clk), .rst(rst), .POP(wire_31), .PUSH(wire_30), .VALUE(wire_3), .OUTPUT(wire_38));
  LEG_ALU # (.UUID(64'd371511248517226547 ^ UUID)) LEG_ALU_68 (.clk(clk), .rst(rst), .\�_____ (wire_58), .\�______1 (wire_0), .\�______2 (wire_10), .Output(wire_111));
  TC_Mux # (.UUID(64'd1931678000695181394 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_69 (.sel(wire_106), .in0(wire_19[7:0]), .in1(wire_2), .out(wire_91));
  TC_And # (.UUID(64'd3760844764780914281 ^ UUID), .BIT_WIDTH(64'd1)) And_70 (.in0(wire_13), .in1(wire_7), .out(wire_106));
  TC_Not # (.UUID(64'd327435945158429862 ^ UUID), .BIT_WIDTH(64'd1)) Not_71 (.in(wire_22), .out(wire_7));
  TC_Equal # (.UUID(64'd3159679139304052043 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_72 (.in0(wire_29), .in1(wire_55), .out(wire_22));
  TC_Equal # (.UUID(64'd1563460054547030821 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_73 (.in0(wire_63), .in1(wire_76), .out(wire_13));
  TC_Splitter8 # (.UUID(64'd1889030559378403173 ^ UUID)) Splitter8_74 (.in(wire_19[7:0]), .out0(wire_112), .out1(wire_100), .out2(wire_99), .out3(wire_101), .out4(), .out5(), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd2004118874441421282 ^ UUID)) Maker8_75 (.in0(wire_112), .in1(wire_100), .in2(wire_99), .in3(wire_101), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_63));
  TC_Splitter8 # (.UUID(64'd1650196065356037064 ^ UUID)) Splitter8_76 (.in(wire_19[7:0]), .out0(), .out1(), .out2(), .out3(), .out4(wire_37), .out5(wire_72), .out6(wire_110), .out7(wire_43));
  TC_Maker8 # (.UUID(64'd4386222698885731789 ^ UUID)) Maker8_77 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(wire_37), .in5(wire_72), .in6(wire_110), .in7(wire_43), .out(wire_29));
  TC_Constant # (.UUID(64'd75759229762736222 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_78 (.out(wire_76));
  TC_Constant # (.UUID(64'd4143237407914741609 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_79 (.out(wire_55));
  TC_Constant # (.UUID(64'd3737133819320673921 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_80 (.out(wire_2));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  wire [7:0] wire_0_4;
  wire [7:0] wire_0_5;
  wire [7:0] wire_0_6;
  wire [7:0] wire_0_7;
  wire [7:0] wire_0_8;
  wire [7:0] wire_0_9;
  wire [7:0] wire_0_10;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6|wire_0_7|wire_0_8|wire_0_9|wire_0_10;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  assign wire_3 = wire_3_0|wire_3_1;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [63:0] wire_8;
  wire [0:0] wire_9;
  assign arch_output_enable = wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_10_0;
  wire [7:0] wire_10_1;
  wire [7:0] wire_10_2;
  wire [7:0] wire_10_3;
  wire [7:0] wire_10_4;
  wire [7:0] wire_10_5;
  wire [7:0] wire_10_6;
  wire [7:0] wire_10_7;
  wire [7:0] wire_10_8;
  wire [7:0] wire_10_9;
  wire [7:0] wire_10_10;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2|wire_10_3|wire_10_4|wire_10_5|wire_10_6|wire_10_7|wire_10_8|wire_10_9|wire_10_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [7:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [63:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [7:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [63:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [7:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [7:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  assign arch_input_enable = wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [7:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [7:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;

endmodule
