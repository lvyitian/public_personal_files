module OVERTUREz_2 (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_24), .en(wire_43), .out(arch_output_value));
  TC_Switch # (.UUID(64'd3 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_33), .in(arch_input_value), .out(wire_26));
  TC_Decoder3 # (.UUID(64'd4053305677990891180 ^ UUID)) Decoder3_2 (.dis(wire_20), .sel0(wire_22), .sel1(wire_12), .sel2(wire_9), .out0(wire_1), .out1(wire_0), .out2(wire_37), .out3(wire_42), .out4(wire_18), .out5(wire_3), .out6(wire_43), .out7());
  TC_Decoder3 # (.UUID(64'd2939524096225771694 ^ UUID)) Decoder3_3 (.dis(wire_20), .sel0(wire_16), .sel1(wire_27), .sel2(wire_4), .out0(wire_45), .out1(wire_51), .out2(wire_50), .out3(wire_23), .out4(wire_41), .out5(wire_30), .out6(wire_33), .out7());
  TC_Splitter8 # (.UUID(64'd1320618894737551008 ^ UUID)) Splitter8_4 (.in(wire_28), .out0(wire_22), .out1(wire_12), .out2(wire_9), .out3(wire_16), .out4(wire_27), .out5(wire_4), .out6(wire_48), .out7(wire_44));
  TC_Maker8 # (.UUID(64'd3189586602702497120 ^ UUID)) Maker8_5 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(wire_48), .in7(wire_44), .out(wire_39));
  TC_Not # (.UUID(64'd478618607012236654 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_47), .out(wire_20));
  TC_Maker8 # (.UUID(64'd3043043946245769206 ^ UUID)) Maker8_7 (.in0(wire_22), .in1(wire_12), .in2(wire_9), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_17));
  TC_Or # (.UUID(64'd3022418375166233711 ^ UUID), .BIT_WIDTH(64'd1)) Or_8 (.in0(wire_42), .in1(wire_13), .out(wire_29));
  TC_Mux # (.UUID(64'd1099724461993398806 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_9 (.sel(wire_13), .in0(wire_24), .in1(wire_40), .out(wire_34));
  TC_Counter # (.UUID(64'd2660306455988799907 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_10 (.clk(clk), .rst(rst), .save(wire_46), .in(wire_31), .out(wire_10));
  TC_Switch # (.UUID(64'd981655355602569219 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(1'd0), .in(1'd0), .out());
  TC_Maker8 # (.UUID(64'd206178571958271433 ^ UUID)) Maker8_12 (.in0(wire_22), .in1(wire_12), .in2(wire_9), .in3(wire_16), .in4(wire_27), .in5(wire_4), .in6(1'd0), .in7(1'd0), .out(wire_5));
  TC_Switch # (.UUID(64'd2794610099783483379 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_36), .in(wire_5), .out(wire_7));
  TC_Mux # (.UUID(64'd3832429127902270701 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_14 (.sel(wire_36), .in0(wire_26), .in1(wire_7), .out(wire_38));
  TC_Or # (.UUID(64'd3773992369932122270 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_1), .in1(wire_36), .out(wire_49));
  TC_Or # (.UUID(64'd1707779249134613013 ^ UUID), .BIT_WIDTH(64'd8)) Or8_16 (.in0(wire_2), .in1(wire_38), .out(wire_24));
  TC_Switch # (.UUID(64'd4288093911554738123 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_11), .in(wire_19), .out(wire_32));
  TC_Not # (.UUID(64'd1174717356322787613 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_11), .out(wire_21));
  TC_Maker8 # (.UUID(64'd1571914357012295039 ^ UUID)) Maker8_19 (.in0(wire_22), .in1(wire_12), .in2(wire_9), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_15));
  TC_Not # (.UUID(64'd2890865550521959735 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_8), .out(wire_14));
  TC_And # (.UUID(64'd2963401396771204859 ^ UUID), .BIT_WIDTH(64'd1)) And_21 (.in0(wire_14), .in1(wire_32), .out(wire_46));
  TC_Decoder3 # (.UUID(64'd3759771637714616433 ^ UUID)) Decoder3_22 (.dis(wire_21), .sel0(wire_22), .sel1(wire_12), .sel2(wire_9), .out0(wire_8), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Program8_1 # (.UUID(64'd5 ^ UUID), .DEFAULT_FILE_NAME("Program8_1_5.w8.bin"), .ARG_SIG("Program8_1_5=%s")) Program8_1_23 (.clk(clk), .rst(rst), .address(wire_10), .out(wire_28));
  DEC # (.UUID(64'd2786871522687439001 ^ UUID)) DEC_24 (.clk(clk), .rst(rst), .OPCODE(wire_39), .IMMEDIATE(wire_36), .CALCULATION(wire_13), .COPY(wire_47), .CONDITION(wire_11));
  ALU # (.UUID(64'd4394841055274257672 ^ UUID)) ALU_25 (.clk(clk), .rst(rst), .\�_____ (wire_17), .\�______1 (wire_6), .\�______2 (wire_25), .Output(wire_40));
  COND # (.UUID(64'd3513967635086646434 ^ UUID)) COND_26 (.clk(clk), .rst(rst), .\�_____ (wire_15), .\�______1 (wire_35), .\�______2 (wire_19));
  RegisterPlus # (.UUID(64'd100000 ^ UUID)) RegisterPlus_27 (.clk(clk), .rst(rst), .\�_____ (wire_45), .\�___________ (wire_24), .\�_____ (wire_49), .\�___________ (wire_31), .Output(wire_2_0));
  RegisterPlus # (.UUID(64'd110000 ^ UUID)) RegisterPlus_28 (.clk(clk), .rst(rst), .\�_____ (wire_51), .\�___________ (wire_24), .\�_____ (wire_0), .\�___________ (wire_6), .Output(wire_2_1));
  RegisterPlus # (.UUID(64'd120000 ^ UUID)) RegisterPlus_29 (.clk(clk), .rst(rst), .\�_____ (wire_50), .\�___________ (wire_24), .\�_____ (wire_37), .\�___________ (wire_25), .Output(wire_2_2));
  RegisterPlus # (.UUID(64'd130000 ^ UUID)) RegisterPlus_30 (.clk(clk), .rst(rst), .\�_____ (wire_23), .\�___________ (wire_34), .\�_____ (wire_29), .\�___________ (wire_35), .Output(wire_2_3));
  RegisterPlus # (.UUID(64'd140000 ^ UUID)) RegisterPlus_31 (.clk(clk), .rst(rst), .\�_____ (wire_41), .\�___________ (wire_24), .\�_____ (wire_18), .\�___________ (), .Output(wire_2_4));
  RegisterPlus # (.UUID(64'd150000 ^ UUID)) RegisterPlus_32 (.clk(clk), .rst(rst), .\�_____ (wire_30), .\�___________ (wire_24), .\�_____ (wire_3), .\�___________ (), .Output(wire_2_5));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  assign arch_input_enable = wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  assign arch_output_enable = wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;

endmodule
