module LEG_COND (clk, rst, ARG1, ARG2, \�_____ , Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] ARG1;
  input  wire [7:0] ARG2;
  input  wire [7:0] \�_____ ;
  output  wire [0:0] Output;

  TC_Equal # (.UUID(64'd469022450449281397 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_0 (.in0(wire_0), .in1(wire_26), .out(wire_27));
  TC_Constant # (.UUID(64'd2051448023974927123 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h20)) Constant8_1 (.out(wire_26));
  TC_Equal # (.UUID(64'd302087503831493541 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_2 (.in0(wire_0), .in1(wire_19), .out(wire_24));
  TC_Constant # (.UUID(64'd4542222613295176889 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h21)) Constant8_3 (.out(wire_19));
  TC_Equal # (.UUID(64'd3977699302148921626 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_4 (.in0(wire_0), .in1(wire_7), .out(wire_4));
  TC_Constant # (.UUID(64'd2314937324333883295 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h22)) Constant8_5 (.out(wire_7));
  TC_Equal # (.UUID(64'd2598179579939704549 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_6 (.in0(wire_0), .in1(wire_18), .out(wire_22));
  TC_Constant # (.UUID(64'd2619140119885518802 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h23)) Constant8_7 (.out(wire_18));
  TC_Equal # (.UUID(64'd1016355148453492596 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_8 (.in0(wire_0), .in1(wire_15), .out(wire_13));
  TC_Constant # (.UUID(64'd1550705849817143486 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h24)) Constant8_9 (.out(wire_15));
  TC_Equal # (.UUID(64'd1602625343120996724 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_10 (.in0(wire_0), .in1(wire_9), .out(wire_8));
  TC_Constant # (.UUID(64'd2222307270319111175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h25)) Constant8_11 (.out(wire_9));
  TC_Not # (.UUID(64'd2244182005895984404 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_12), .out(wire_23));
  TC_Equal # (.UUID(64'd168532653866922664 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_13 (.in0(wire_14), .in1(wire_1), .out(wire_12));
  TC_Switch # (.UUID(64'd859839441511864255 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_27), .in(wire_12), .out(wire_5_0));
  TC_Switch # (.UUID(64'd3687602544865986092 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_15 (.en(wire_24), .in(wire_23), .out(wire_5_1));
  TC_LessU # (.UUID(64'd2837489368470343284 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_16 (.in0(wire_14), .in1(wire_1), .out(wire_2));
  TC_Switch # (.UUID(64'd114564404545293814 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_4), .in(wire_2), .out(wire_5_2));
  TC_Switch # (.UUID(64'd3233876504730006742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_22), .in(wire_17), .out(wire_5_5));
  TC_Or # (.UUID(64'd1752390656836275508 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_2), .in1(wire_12), .out(wire_17));
  TC_Switch # (.UUID(64'd1313143816079393951 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_20 (.en(wire_8), .in(wire_3), .out(wire_5_3));
  TC_Not # (.UUID(64'd1225463839904331438 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_2), .out(wire_3));
  TC_Switch # (.UUID(64'd3591175240098488323 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_13), .in(wire_16), .out(wire_5_4));
  TC_And # (.UUID(64'd2923998825401666618 ^ UUID), .BIT_WIDTH(64'd1)) And_23 (.in0(wire_23), .in1(wire_3), .out(wire_16));
  TC_Maker8 # (.UUID(64'd4350048876850400171 ^ UUID)) Maker8_24 (.in0(wire_21), .in1(wire_28), .in2(wire_6), .in3(wire_20), .in4(wire_10), .in5(wire_11), .in6(1'd0), .in7(1'd0), .out(wire_0));
  TC_Splitter8 # (.UUID(64'd3964202440971776894 ^ UUID)) Splitter8_25 (.in(wire_25), .out0(wire_21), .out1(wire_28), .out2(wire_6), .out3(wire_20), .out4(wire_10), .out5(wire_11), .out6(), .out7());

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  assign wire_1 = ARG2;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_5_0;
  wire [0:0] wire_5_1;
  wire [0:0] wire_5_2;
  wire [0:0] wire_5_3;
  wire [0:0] wire_5_4;
  wire [0:0] wire_5_5;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3|wire_5_4|wire_5_5;
  assign Output = wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  assign wire_14 = ARG1;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  assign wire_25 = \�_____ ;
  wire [7:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;

endmodule
