module LEG_COND (clk, rst, ARG1, ARG2, \�_____ , Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] ARG1;
  input  wire [7:0] ARG2;
  input  wire [7:0] \�_____ ;
  output  wire [0:0] Output;

  TC_Equal # (.UUID(64'd469022450449281397 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_0 (.in0(wire_3), .in1(wire_20), .out(wire_15));
  TC_Constant # (.UUID(64'd2051448023974927123 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h20)) Constant8_1 (.out(wire_20));
  TC_Equal # (.UUID(64'd302087503831493541 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_2 (.in0(wire_3), .in1(wire_13), .out(wire_5));
  TC_Constant # (.UUID(64'd4542222613295176889 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h21)) Constant8_3 (.out(wire_13));
  TC_Equal # (.UUID(64'd3977699302148921626 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_4 (.in0(wire_3), .in1(wire_17), .out(wire_7));
  TC_Constant # (.UUID(64'd2314937324333883295 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h22)) Constant8_5 (.out(wire_17));
  TC_Equal # (.UUID(64'd2598179579939704549 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_6 (.in0(wire_3), .in1(wire_19), .out(wire_12));
  TC_Constant # (.UUID(64'd2619140119885518802 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h23)) Constant8_7 (.out(wire_19));
  TC_Equal # (.UUID(64'd1016355148453492596 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_8 (.in0(wire_3), .in1(wire_4), .out(wire_14));
  TC_Constant # (.UUID(64'd1550705849817143486 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h24)) Constant8_9 (.out(wire_4));
  TC_Equal # (.UUID(64'd1602625343120996724 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_10 (.in0(wire_3), .in1(wire_10), .out(wire_9));
  TC_Constant # (.UUID(64'd2222307270319111175 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h25)) Constant8_11 (.out(wire_10));
  TC_Not # (.UUID(64'd2244182005895984404 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_1), .out(wire_21));
  TC_Equal # (.UUID(64'd168532653866922664 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_13 (.in0(wire_0), .in1(wire_8), .out(wire_1));
  TC_Switch # (.UUID(64'd859839441511864255 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_15), .in(wire_1), .out(wire_6_0));
  TC_Switch # (.UUID(64'd3687602544865986092 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_15 (.en(wire_5), .in(wire_21), .out(wire_6_4));
  TC_LessU # (.UUID(64'd2837489368470343284 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_16 (.in0(wire_0), .in1(wire_8), .out(wire_2));
  TC_Switch # (.UUID(64'd114564404545293814 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_7), .in(wire_2), .out(wire_6_5));
  TC_Switch # (.UUID(64'd3233876504730006742 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_12), .in(wire_16), .out(wire_6_3));
  TC_Or # (.UUID(64'd1752390656836275508 ^ UUID), .BIT_WIDTH(64'd1)) Or_19 (.in0(wire_2), .in1(wire_1), .out(wire_16));
  TC_Switch # (.UUID(64'd1313143816079393951 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_20 (.en(wire_9), .in(wire_18), .out(wire_6_1));
  TC_Not # (.UUID(64'd1225463839904331438 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_2), .out(wire_18));
  TC_Switch # (.UUID(64'd3591175240098488323 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_14), .in(wire_11), .out(wire_6_2));
  TC_And # (.UUID(64'd2923998825401666618 ^ UUID), .BIT_WIDTH(64'd1)) And_23 (.in0(wire_21), .in1(wire_18), .out(wire_11));

  wire [7:0] wire_0;
  assign wire_0 = ARG1;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  assign wire_3 = \�_____ ;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_6_0;
  wire [0:0] wire_6_1;
  wire [0:0] wire_6_2;
  wire [0:0] wire_6_3;
  wire [0:0] wire_6_4;
  wire [0:0] wire_6_5;
  assign wire_6 = wire_6_0|wire_6_1|wire_6_2|wire_6_3|wire_6_4|wire_6_5;
  assign Output = wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  assign wire_8 = ARG2;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;

endmodule
