module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_20), .en(wire_53), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_110), .in(arch_input_value), .out(wire_116));
  TC_Counter # (.UUID(64'd1175999672554394000 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_2 (.clk(clk), .rst(rst), .save(wire_9), .in(wire_20), .out(wire_24));
  TC_Splitter8 # (.UUID(64'd3496280010280654809 ^ UUID)) Splitter8_3 (.in(wire_12), .out0(wire_4), .out1(wire_67), .out2(wire_38), .out3(wire_101), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1350359362790102949 ^ UUID)) Splitter8_4 (.in(wire_33), .out0(wire_78), .out1(wire_72), .out2(wire_112), .out3(wire_63), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3688384451292696869 ^ UUID)) Splitter8_5 (.in(wire_117), .out0(wire_15), .out1(wire_99), .out2(wire_30), .out3(wire_88), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3357720912797461292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_61), .in(wire_24), .out());
  TC_Maker8 # (.UUID(64'd2922775923237819214 ^ UUID)) Maker8_7 (.in0(wire_106), .in1(wire_81), .in2(wire_50), .in3(wire_49), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_1));
  TC_Splitter8 # (.UUID(64'd4136660363423911410 ^ UUID)) Splitter8_8 (.in(wire_77[7:0]), .out0(wire_106), .out1(wire_81), .out2(wire_50), .out3(wire_49), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd4550958897663313502 ^ UUID)) Splitter8_9 (.in(wire_77[7:0]), .out0(wire_71), .out1(wire_69), .out2(wire_103), .out3(wire_42), .out4(wire_46), .out5(wire_57), .out6(wire_65), .out7(wire_14));
  TC_Maker8 # (.UUID(64'd3153840370766490713 ^ UUID)) Maker8_10 (.in0(wire_71), .in1(wire_69), .in2(wire_103), .in3(wire_42), .in4(wire_46), .in5(wire_57), .in6(wire_65), .in7(wire_14), .out(wire_92));
  TC_Constant # (.UUID(64'd4029987529778329422 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out(wire_16));
  TC_Constant # (.UUID(64'd47372170638122597 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out(wire_105));
  TC_Constant # (.UUID(64'd3010400910295959985 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_19));
  TC_Constant # (.UUID(64'd1353887318054096472 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_7));
  TC_Constant # (.UUID(64'd4461919415197064488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out(wire_74));
  TC_Constant # (.UUID(64'd2551986311311524963 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_37));
  TC_Switch # (.UUID(64'd201407107924193690 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_102), .in(wire_40), .out(wire_28_0));
  TC_Switch # (.UUID(64'd3784926049681585699 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_93), .in(wire_40), .out(wire_3_0));
  TC_Switch # (.UUID(64'd3418942253385023549 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_10), .in(wire_86), .out(wire_28_5));
  TC_Switch # (.UUID(64'd3104771108315787100 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_6), .in(wire_86), .out(wire_3_10));
  TC_Switch # (.UUID(64'd494263610589549334 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_121), .in(wire_76), .out(wire_28_6));
  TC_Switch # (.UUID(64'd4455028313033582898 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_64), .in(wire_76), .out(wire_3_6));
  TC_Switch # (.UUID(64'd977062972681925203 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_35), .in(wire_31), .out(wire_28_8));
  TC_Switch # (.UUID(64'd2935373336597064260 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_119), .in(wire_31), .out(wire_3_9));
  TC_Switch # (.UUID(64'd2595310988575568445 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_13), .in(wire_91), .out(wire_28_7));
  TC_Switch # (.UUID(64'd3649926646471230167 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_56), .in(wire_91), .out(wire_3_8));
  TC_Switch # (.UUID(64'd115863760055946247 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_80), .in(wire_26), .out(wire_28_9));
  TC_Switch # (.UUID(64'd459043271910661458 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_5), .in(wire_26), .out(wire_3_7));
  TC_Switch # (.UUID(64'd4275937720180353902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_66), .in(wire_24), .out());
  TC_Switch # (.UUID(64'd2718446434835356700 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_27), .in(wire_116), .out(wire_28_10));
  TC_Switch # (.UUID(64'd1811299859375739998 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_84), .in(wire_116), .out(wire_3_5));
  TC_Or # (.UUID(64'd117421755651659184 ^ UUID), .BIT_WIDTH(64'd1)) Or_32 (.in0(wire_27), .in1(wire_84), .out(wire_110));
  TC_Switch # (.UUID(64'd262409980643160938 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_36), .in(wire_34[7:0]), .out(wire_3_3));
  TC_Switch # (.UUID(64'd2764614579549035605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_48), .in(wire_58[7:0]), .out(wire_28_1));
  TC_Switch # (.UUID(64'd2974460371787013801 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_45), .in(wire_118), .out(wire_20_0));
  TC_Mux # (.UUID(64'd1769789085559769130 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_36 (.sel(wire_36), .in0(wire_34[7:0]), .in1(wire_59), .out(wire_33));
  TC_Mux # (.UUID(64'd1404337327044278632 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_37 (.sel(wire_48), .in0(wire_58[7:0]), .in1(wire_0), .out(wire_12));
  TC_Constant # (.UUID(64'd4387708643330744374 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_38 (.out(wire_0));
  TC_Constant # (.UUID(64'd2430039925245603401 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_39 (.out(wire_59));
  TC_Switch # (.UUID(64'd3877536405880520929 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_29), .in(wire_120), .out(wire_23));
  TC_Constant # (.UUID(64'd2430392602802046886 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_41 (.out(wire_18));
  TC_Mux # (.UUID(64'd1559488034901936773 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_42 (.sel(wire_23), .in0(wire_52), .in1(wire_18), .out(wire_117));
  TC_Switch # (.UUID(64'd3981948550050450551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_23), .in(wire_25[7:0]), .out(wire_20_1));
  TC_Ram # (.UUID(64'd1683242105781375453 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_44 (.clk(clk), .rst(rst), .load(wire_43), .save(wire_62), .address({{24{1'b0}}, wire_104 }), .in0({{56{1'b0}}, wire_20 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_95), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd1949247607308932292 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_45 (.out(wire_111));
  TC_Or # (.UUID(64'd2571069615494455195 ^ UUID), .BIT_WIDTH(64'd1)) Or_46 (.in0(wire_41), .in1(wire_22), .out(wire_43));
  TC_Switch # (.UUID(64'd3896516251333244950 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_73), .in(wire_11), .out(wire_28_4));
  TC_Switch # (.UUID(64'd4219278115069450234 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_100), .in(wire_11), .out(wire_3_1));
  TC_Switch # (.UUID(64'd875265095609107539 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_41), .in(wire_95[7:0]), .out(wire_28_3));
  TC_Switch # (.UUID(64'd1025433274855748469 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_22), .in(wire_95[7:0]), .out(wire_3_4));
  TC_Program # (.UUID(64'd4489305393227859486 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_3E4D37784397861E.w8.bin"), .ARG_SIG("Program_3E4D37784397861E=%s")) Program_51 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_24 }), .out0(wire_77), .out1(wire_58), .out2(wire_34), .out3(wire_25));
  TC_Switch # (.UUID(64'd3036050060892365836 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_54), .in(wire_44), .out(wire_28_2));
  TC_Switch # (.UUID(64'd3830579770898048556 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_2), .in(wire_44), .out(wire_3_2));
  TC_Or # (.UUID(64'd1511395350716789461 ^ UUID), .BIT_WIDTH(64'd1)) Or_54 (.in0(wire_54), .in1(wire_2), .out(wire_98));
  TC_Mux # (.UUID(64'd1931678000695181394 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_55 (.sel(wire_97), .in0(wire_25[7:0]), .in1(wire_114), .out(wire_52));
  TC_And # (.UUID(64'd3760844764780914281 ^ UUID), .BIT_WIDTH(64'd1)) And_56 (.in0(wire_21), .in1(wire_39), .out(wire_60));
  TC_Not # (.UUID(64'd327435945158429862 ^ UUID), .BIT_WIDTH(64'd1)) Not_57 (.in(wire_113), .out(wire_39));
  TC_Equal # (.UUID(64'd3159679139304052043 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_58 (.in0(wire_47), .in1(wire_55), .out(wire_113));
  TC_Equal # (.UUID(64'd1563460054547030821 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_59 (.in0(wire_87), .in1(wire_85), .out(wire_21));
  TC_Splitter8 # (.UUID(64'd1889030559378403173 ^ UUID)) Splitter8_60 (.in(wire_25[7:0]), .out0(wire_51), .out1(wire_115), .out2(wire_107), .out3(wire_83), .out4(), .out5(), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd2004118874441421282 ^ UUID)) Maker8_61 (.in0(wire_51), .in1(wire_115), .in2(wire_107), .in3(wire_83), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_87));
  TC_Splitter8 # (.UUID(64'd1650196065356037064 ^ UUID)) Splitter8_62 (.in(wire_25[7:0]), .out0(), .out1(), .out2(), .out3(), .out4(wire_94), .out5(wire_75), .out6(wire_108), .out7(wire_17));
  TC_Maker8 # (.UUID(64'd4386222698885731789 ^ UUID)) Maker8_63 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(wire_94), .in5(wire_75), .in6(wire_108), .in7(wire_17), .out(wire_47));
  TC_Constant # (.UUID(64'd75759229762736222 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_64 (.out(wire_85));
  TC_Constant # (.UUID(64'd4143237407914741609 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_65 (.out(wire_55));
  TC_Constant # (.UUID(64'd3737133819320673921 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hF)) Constant8_66 (.out(wire_114));
  TC_Or # (.UUID(64'd1560433342647392432 ^ UUID), .BIT_WIDTH(64'd1)) Or_67 (.in0(wire_79), .in1(wire_60), .out(wire_97));
  TC_And # (.UUID(64'd2200126785490710302 ^ UUID), .BIT_WIDTH(64'd1)) And_68 (.in0(wire_70), .in1(wire_29), .out(wire_79));
  TC_Not # (.UUID(64'd1299938039481718942 ^ UUID), .BIT_WIDTH(64'd1)) Not_69 (.in(wire_23), .out(wire_70));
  _4bit_Decoder # (.UUID(64'd188593635878702660 ^ UUID)) _4bit_Decoder_70 (.clk(clk), .rst(rst), .\1_1 (wire_4), .\2_1 (wire_67), .\4_1 (wire_38), .\8_1 (wire_101), .\7 (wire_27), .\11 (), .\3 (wire_35), .\15 (), .\6 (wire_61), .\8_2 (wire_73), .\5 (wire_80), .\9 (wire_41), .\10 (wire_54), .\4_2 (wire_13), .\12 (), .\13 (), .\14 (), .\2_2 (wire_121), .\1_2 (wire_10), .\0 (wire_102));
  _4bit_Decoder # (.UUID(64'd3657203059375966986 ^ UUID)) _4bit_Decoder_71 (.clk(clk), .rst(rst), .\1_1 (wire_78), .\2_1 (wire_72), .\4_1 (wire_112), .\8_1 (wire_63), .\7 (wire_84), .\11 (), .\3 (wire_119), .\15 (), .\6 (wire_66), .\8_2 (wire_100), .\5 (wire_5), .\9 (wire_22), .\10 (wire_2), .\4_2 (wire_56), .\12 (), .\13 (), .\14 (), .\2_2 (wire_64), .\1_2 (wire_6), .\0 (wire_93));
  _4bit_Decoder # (.UUID(64'd4526675728054865805 ^ UUID)) _4bit_Decoder_72 (.clk(clk), .rst(rst), .\1_1 (wire_15), .\2_1 (wire_99), .\4_1 (wire_30), .\8_1 (wire_88), .\7 (wire_53), .\11 (), .\3 (wire_32), .\15 (), .\6 (wire_9), .\8_2 (wire_90), .\5 (wire_8), .\9 (wire_62), .\10 (wire_96), .\4_2 (wire_82), .\12 (), .\13 (), .\14 (), .\2_2 (wire_68), .\1_2 (wire_89), .\0 (wire_109));
  RegisterPlus # (.UUID(64'd1898575026262245003 ^ UUID)) RegisterPlus_73 (.clk(clk), .rst(rst), .\�_____ (wire_16), .\�___________ (wire_20), .\�_____ (wire_109), .\�___________ (), .Output(wire_40));
  RegisterPlus # (.UUID(64'd201486149512558618 ^ UUID)) RegisterPlus_74 (.clk(clk), .rst(rst), .\�_____ (wire_105), .\�___________ (wire_20), .\�_____ (wire_89), .\�___________ (), .Output(wire_86));
  RegisterPlus # (.UUID(64'd4130910523704063521 ^ UUID)) RegisterPlus_75 (.clk(clk), .rst(rst), .\�_____ (wire_19), .\�___________ (wire_20), .\�_____ (wire_68), .\�___________ (), .Output(wire_76));
  RegisterPlus # (.UUID(64'd579904311903668382 ^ UUID)) RegisterPlus_76 (.clk(clk), .rst(rst), .\�_____ (wire_7), .\�___________ (wire_20), .\�_____ (wire_32), .\�___________ (), .Output(wire_31));
  RegisterPlus # (.UUID(64'd2026589517635316452 ^ UUID)) RegisterPlus_77 (.clk(clk), .rst(rst), .\�_____ (wire_74), .\�___________ (wire_20), .\�_____ (wire_82), .\�___________ (), .Output(wire_91));
  RegisterPlus # (.UUID(64'd1622410096212380183 ^ UUID)) RegisterPlus_78 (.clk(clk), .rst(rst), .\�_____ (wire_37), .\�___________ (wire_20), .\�_____ (wire_8), .\�___________ (), .Output(wire_26));
  LEG_COND # (.UUID(64'd999600516743479399 ^ UUID)) LEG_COND_79 (.clk(clk), .rst(rst), .ARG1(wire_28), .ARG2(wire_3), .\�_____ (wire_77[7:0]), .Output(wire_120));
  RegisterPlus # (.UUID(64'd471658098348471390 ^ UUID)) RegisterPlus_80 (.clk(clk), .rst(rst), .\�_____ (wire_111), .\�___________ (wire_20), .\�_____ (wire_90), .\�___________ (wire_104), .Output(wire_11));
  LEG_DEC # (.UUID(64'd2015393024950033718 ^ UUID)) LEG_DEC_81 (.clk(clk), .rst(rst), .OPCODE(wire_92), .IMMEDIATE1(wire_48), .IMMEDIATE2(wire_36), .CALCULATION(wire_45), .JUMP(wire_29));
  LEG_ALU # (.UUID(64'd371511248517226547 ^ UUID)) LEG_ALU_82 (.clk(clk), .rst(rst), .\�_____ (wire_1), .\�______1 (wire_28), .\�______2 (wire_3), .Output(wire_118));
  ZXE6ZXA0ZX88 # (.UUID(64'd1554391434741513408 ^ UUID)) ZXE6ZXA0ZX88_83 (.clk(clk), .rst(rst), .POP(wire_98), .PUSH(wire_96), .VALUE(wire_20), .OUTPUT(wire_44));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  wire [7:0] wire_3_8;
  wire [7:0] wire_3_9;
  wire [7:0] wire_3_10;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7|wire_3_8|wire_3_9|wire_3_10;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_20_0;
  wire [7:0] wire_20_1;
  assign wire_20 = wire_20_0|wire_20_1;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [63:0] wire_25;
  wire [7:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_28_0;
  wire [7:0] wire_28_1;
  wire [7:0] wire_28_2;
  wire [7:0] wire_28_3;
  wire [7:0] wire_28_4;
  wire [7:0] wire_28_5;
  wire [7:0] wire_28_6;
  wire [7:0] wire_28_7;
  wire [7:0] wire_28_8;
  wire [7:0] wire_28_9;
  wire [7:0] wire_28_10;
  assign wire_28 = wire_28_0|wire_28_1|wire_28_2|wire_28_3|wire_28_4|wire_28_5|wire_28_6|wire_28_7|wire_28_8|wire_28_9|wire_28_10;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [63:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  assign arch_output_enable = wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [63:0] wire_58;
  wire [7:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [7:0] wire_76;
  wire [63:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [7:0] wire_85;
  wire [7:0] wire_86;
  wire [7:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;
  wire [7:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [63:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [7:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  assign arch_input_enable = wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [7:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [7:0] wire_117;
  wire [7:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;

endmodule
