module LEG_DEC (clk, rst, OPCODE, IMMEDIATE1, IMMEDIATE2, CALCULATION, JUMP);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] OPCODE;
  output  wire [0:0] IMMEDIATE1;
  output  wire [0:0] IMMEDIATE2;
  output  wire [0:0] CALCULATION;
  output  wire [0:0] JUMP;

  TC_Splitter8 # (.UUID(64'd2459092867252704659 ^ UUID)) Splitter8_0 (.in(wire_25), .out0(), .out1(), .out2(), .out3(), .out4(wire_3), .out5(wire_2), .out6(wire_20), .out7(wire_0));
  TC_Equal # (.UUID(64'd4451411414923206213 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_1 (.in0(wire_1), .in1(wire_24), .out(wire_13));
  TC_Constant # (.UUID(64'd4146811536148831861 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h20)) Constant8_2 (.out(wire_24));
  TC_Equal # (.UUID(64'd3175768114047069080 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_3 (.in0(wire_1), .in1(wire_10), .out(wire_27));
  TC_Constant # (.UUID(64'd2100458896617105062 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h21)) Constant8_4 (.out(wire_10));
  TC_Equal # (.UUID(64'd18612831955176227 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_5 (.in0(wire_1), .in1(wire_26), .out(wire_22));
  TC_Constant # (.UUID(64'd4436786725961600454 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h22)) Constant8_6 (.out(wire_26));
  TC_Equal # (.UUID(64'd3951549131992813285 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_7 (.in0(wire_1), .in1(wire_16), .out(wire_9));
  TC_Constant # (.UUID(64'd2187694636879553517 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h23)) Constant8_8 (.out(wire_16));
  TC_Equal # (.UUID(64'd1722280921780021930 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_9 (.in0(wire_1), .in1(wire_7), .out(wire_12));
  TC_Constant # (.UUID(64'd1232993965608782474 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h24)) Constant8_10 (.out(wire_7));
  TC_Equal # (.UUID(64'd1677764983551709104 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_11 (.in0(wire_1), .in1(wire_14), .out(wire_23));
  TC_Constant # (.UUID(64'd3969712149290372119 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h25)) Constant8_12 (.out(wire_14));
  TC_Or3 # (.UUID(64'd4231655371929136514 ^ UUID), .BIT_WIDTH(64'd1)) Or3_13 (.in0(wire_13), .in1(wire_27), .in2(wire_22), .out(wire_18));
  TC_Or3 # (.UUID(64'd493742362470177643 ^ UUID), .BIT_WIDTH(64'd1)) Or3_14 (.in0(wire_18), .in1(wire_9), .in2(wire_12), .out(wire_5));
  TC_Or # (.UUID(64'd3897193912910816394 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_5), .in1(wire_23), .out(wire_19));
  _4bit_Decoder # (.UUID(64'd2481737798594514154 ^ UUID)) _4bit_Decoder_16 (.clk(clk), .rst(rst), .\1_1 (wire_3), .\2_1 (wire_2), .\4_1 (1'd0), .\8_1 (1'd0), .\7 (), .\11 (), .\3 (), .\15 (), .\6 (), .\8_2 (), .\5 (), .\9 (), .\10 (), .\4_2 (), .\12 (), .\13 (), .\14 (), .\2_2 (), .\1_2 (), .\0 (wire_4));
  TC_Maker8 # (.UUID(64'd2291807996615366193 ^ UUID)) Maker8_17 (.in0(wire_15), .in1(wire_21), .in2(wire_11), .in3(wire_17), .in4(wire_6), .in5(wire_8), .in6(1'd0), .in7(1'd0), .out(wire_1));
  TC_Splitter8 # (.UUID(64'd4080107753313342668 ^ UUID)) Splitter8_18 (.in(wire_25), .out0(wire_15), .out1(wire_21), .out2(wire_11), .out3(wire_17), .out4(wire_6), .out5(wire_8), .out6(), .out7());

  wire [0:0] wire_0;
  assign IMMEDIATE1 = wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  assign CALCULATION = wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  assign JUMP = wire_19;
  wire [0:0] wire_20;
  assign IMMEDIATE2 = wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  assign wire_25 = OPCODE;
  wire [7:0] wire_26;
  wire [0:0] wire_27;

endmodule
